`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2LeHPrWCYe5+ReQ8YltqsvkIJm1v+VBYBDVzugbhOoXx3pBXXWE4qI6F8fYSidcj
coDVWgRSg1vzUY1OxgD72JoNu5LAe4lBuybfcig2TzY9p/Xx7ohwGhD8dXG7sBaT
Yt2V9V9leDUO5Kfbi/eGMTHewqSbeK5y6VMQzgT+2nu7Pl8+/W+7fQclXeeipdLS
IY2f2mOcHSVGVvsgNOJkSgxvDK7McL6kKSq+a1ezn02PEYBsbBGqcx+KFKO0Fpgl
Z4DKUQmv/isKU6LKq/f3FmOpqYrsbo/spdc/sAD+pRt+MBAcvFKt8Hy3dSWTZfGB
qVU0ZuLCTbYZNSKIHF7x4sLhthznGK/9XVH3rUzwrSVsDNCiJ1IyPqrQYUNbTBXj
cayqESBclXcK6dQokvDpuO0Pa3yCWfFJPehLCkHb9cgbGeA9vdJJKFWg4MxEHvIw
yNBfAG1a6GgCDImlETeuUrYygVZd0quJXdVBUqtasXh9/seeHqLl9+l4lD8ySCUw
sgkheoepHEm8Rd7obeUS/cAWkIcd8Acwo/0FDw6q/JJBWDz5TM9LUOPsP6ISMypB
KzP75YSWSmlUSMzyJ0h9M8CodtJVJh/1zjWaYebt0jh7K0gukcV5MPD7MtIej4aQ
A3qYMmVvFCY70SQVx02QjpuJKKQaNSpb3UMvEK1b+mhuzOJxu2UXF8VmQuO0ER/y
MUW45t0XKp7iIHf3HkOH9YiQ/a67qTwnrQZ8vnsenYDGMH4+5VBbgQCIohuOv3CQ
5xxiE6iQEWOGQOKqFmT+oK/vQjTjm6PSTIHCm3ELE5+ZOLjmw433Ii6+hrUwjaoY
t/msVYEqpwQbCpMMYq4TLtBYM/+q5/5poq+eOtYD5lfXwaumQUm2FMOf3KA3RXaG
Wa8FCJUasIxVpi9ljfzdoNtwcs2VEjWxlTtmw9iDpIoGjKF8kAI4yuLzQsM3gAuc
KPFMf6xhj0H4PyUP9UQ04WHfQmCwetlWKbvXy/WNTuwLk8KIxclPKYxl/u1UqkAl
39mo4Dx5be+QvyE1KZgLu6KUUzZe2RbFgJ5Kl14FmEF1sJ1lFHJplmDsRx9mQgQy
4UTkPRl5WRhARRE7IMzfzWY+KgCSY4xNwEBnjc78FTFpyg3LVxTsWHznuiLpMNlZ
oJzNZu+BaKazNXRTmlIKgilmMDP6nFpY/u0lvbu0lwq1DfWZPbDaiG8GOsT9MqmB
Yxpy/PhvIosTspNG0Zl6IHsY26DnALr5YMndYtZ3NDx9P7RR2FyH7UzeqT8dgIS/
aHMEqxxL3JnpU1gemHXJ3CXxznqPCwBopgVCxUklgmcJl8C8nkS6/vm97Hce3cuJ
rQGcIFa8r5SvATdaxUwEV1TqF3wFd0YCum4kOI94qosjr07Ihwy5JZYpKjuMwDln
1cB0ZhmqPaWHa9u7NV7zfMknaTRF+sGGoHBSFASpABs8JLNwh9WTqL2J7C63DPeY
84zge8dHmP9UUxfCZbTNEXB5LUOhVSSBSTlaBd6XareYR4eb/jYO70JsK9Dst8ao
CcCAdjZ1lHmcgSUXAM03RVNy7VvMZ5IlRq8yXsqu9RL/88Yy31+dBpR9lzY2hxKx
cEiZ9asRvCy99T6GhGcIgLtiNNzq7Aw5QpOnO/l67KVdZvcnINvIhUMvYftSczY5
y+R/XeVqEVFx8PbpK7bF749TMGvo5Eg6Lux7gFaniJgTuYfiuw8rHzobkb5LTta0
7ybIlrVP7XedX0lxN1wUFpfGDIYQyMy3PItTbwSAZp8n9lonQlAYiHFaP2+EIhA1
4TOvwB3rJ8ddiE1IAXaYf2LhqqO8y9ixlLbrjQ6+8vXsHeR3M5WR74WFUgeS7vRR
esbi6jbMj7kmB4Oa/iYvEMTOi8hHpeDf41kWwUg+1NgnnVg5+XWxCfG4pG2zxuLm
rebEfME7L8USmcc0fzyG+c6AjQqhvcJnYkmBWzdHByrW0ykczRoHWA4yLUcsFMK0
4d9VVkeElJUxv4YJqdS9QQ==
`protect END_PROTECTED
