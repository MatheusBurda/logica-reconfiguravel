`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fiePLQNmWaQTeaWv+gK4laJ9uTAI2X047PKy9MB5R+KdMcFqzfI5xUal98as1N0t
YqyDgagwp4TyxYA9w8QULfXK9vCMttedg+VMmIvltCR4/7ZHVR1sqAtDTjwFKTZh
XvThTndvUxhUc5ARgPxD452/GAYM2oWXGViTYLAZPMBz354xD+43318fUgU9RbD6
eQNWa+D3A32UNhWVJw/Pf8LkOrOWKZfIqFZz3BEyYE6JLIN09Ef5Ix99U4hjx5hb
mVML046/5m0oYoNPMI5cNcgsvQLAHuQuSRgbu6VPNmw7G7F4F4pxtPUlbMiwd00Q
litG97vQ5EDok3fHTRJrYo5cOyX2wOWEye+/OBUfindAz3VaHYXcsvVoqM1ij6EM
CtxhGy4dwKILHad4y0HxxF/DgIg9A8nfaoJwqh7RCh7IxOV21mxw7BN+1E2PqgiM
ObywZnSf/zVuU6xi7qPEmj0E4ei5PXWv5wa0Es4to3lfcLm1GAbLoHdI9FAsI4KY
4OJ2ZH2e5OdNlTcyWP8Ea4J2iU9CWAjcDWx4M+mcqrCcah61SIl6L6P8i/SvPXsf
LZy2IbYDH/h/0yvfHt5qqOZKc9FhCDm1vib3MeVrCsktJwJxQG9N2FKckRRqiX7i
JasPfEw+GxgA/uIyOLXnIvwJqextUqZzLz/xgNZLEzkBTEfVXrWDiG4BWolnlqcb
ci+2pDPWyIV6gHALwVAxlhcv9PbRPNT5VolxfEph9H2Laaf3J2BZ5gPJnyQ+i/+b
H9nB55BMMu5US50b6WrkJMSniJiw/y3FG+DtpbJ8JmJrFUxlQzaeyvla9v61frD1
hbpbUUXEUcnTVWuN3FgfKs23yDs+wcoiiI80x3Ceo3LQ5da2cHgDjgJfDP3pQ0BE
IWM3GFaB4a9SttSiPle17O+D2jz54T0m40oFdTRPoR8nx73nxmjZke+MaeylVP4M
s0XJqdFdW+QoPgc+wPKW8TLjTbad00QB/QFUD9TUjohi4puS80H2l6QlWVOnTbEH
y4rDPIyKlL9luviuKWTDUwRQ6gJjt8NLytvufR8BS9wQrA1U4rHIVwVjUar44Not
KO4MYPxBATcj+XA3VpELyvcgmhplCi6jDaWfmzPdTEsl/O4Nw3LoQccgHY/z9Sq9
dGzIj6HlvF1vKtV2jEYn/mGVEMRvjHtRDBa8DWg+EZXaXQB6XxgEO7+FDuocK2Ig
ZEOf/QAikuEA7gXdZw1d+R8oJJAISoqbyCbPN+44Lx7XokqQn6r46vxsHTD4LWGb
pw6ZuKP1LfNXWtXjP4FlZVzBenBM6K5rXTwyP5iOrKs2ZoSxCnRRqusbCdf3zESP
jlpxNkUk2W36nBe8RQ4RykH8s5qdkxy4JOWi3qEoveGSagJPIvSQOg/B6BQIvOvR
AQkeMGCCwDz4suy9Nf5Av0PbsxrS8BPzR2qG/AhIN54vVF7+d3+2C4yDH+x8ZwSe
iiAoAho9psKK0AD8lOMMpxkmmf1lY1qzsVut/ZJ5WTXepb5JJ93oe3nPrrmSCzQ/
d8As4AX83kD7UlsH4zaz1XeprpCwsXEW7S/hwuLyqWnbqyd/Xrrhng+wDDIB10dN
SCVeejhbOjZ0chhQS3jwcWtgI81sWd2GRjmDKnBg7a1jlztCBbjBlQf2L6JRDgLl
pSkmMXyWNHMdvLJ13Lbb034zQWDCVlok5ohUOcMYw8PPuE4kG5V696siekRGIFBm
LDEuJjsp4iyjvD5KFDegzL42mXudRMRWe+zSNxSYFUKEu3VLU8NJsDLwtRT4DQzw
d4U7HeHbTz7tNNjz6PFQdtbiGJg83u66GaRFVHdkQ9BLATy+LvGrniFimapFCKPZ
zkSegC0oj6y5y9S8GXY9lqxAogqf/AC+rhvpXhjC9ktkV6U71DwwFD7QlR0m8cH+
YfzKNRKoKzb63tKU78LMR5ADOalV/l9A6vg92/w/72Yap7Orlaj3BvHIjQh6EBkb
fLPZAjs3cnfBgXjDLFPd6GxXhh5DD9tf3OFqgb03WDW4HaIsSvDfIYlWaflobWJY
5o3hogSoWsoWwu8+PUFwfevl11HXpJn18ODlJnJVQYn2rn/7warzBausK1WNvfL8
T4uKMYSUprJqKWepKw8seXizE7eNyFf12ZhXduUZzlMSh8/SQnIqG7ngRBoQlLAb
4pvz8KavjQmW6UBE8RWQ8XaEbdEjySALgdbo0Ph+XHW8bLfGD4oGBUWNh7Jp1qHF
kGs6rY4ZrZGVaVZr77DhJA==
`protect END_PROTECTED
