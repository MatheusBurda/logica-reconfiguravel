`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n7Ub7JKUKjr3OGo/AhQuPYsIdqX8gnre8RjCmJuZrYbNz0cQOnMnBFK2NCu9DMHo
rQqxMDBp9tnUxNUSAvltMSNA65aee1o7B24N+TRnU4csa3zdO5twUzz6Q9XrRgwF
Yp9+ynYU+DhJ7HYwts/vBOJpzeaxVF/hNGrIp/Qn9O2Y+E5MvgeLsshQHLLcA9NP
h79ut5OY56zIZddJhc4lAqJNmam7H5ku+1v/Lu4eCL97miVt1BR5MNqil7xNDfJh
cHU0auUfBXCjgoJecgrYlwoKsurWYRxEWCbBknJ/vbF4WNgFu/KAPZm4fFdYObP4
rXYr6m/O2GEqrF/7K5wJ87vc6mhqZjOzsbpI01F5HseEm0wvL55kGZtZgjie1BlK
k3s76GMIKHIyWW17ZM92pb5tn2aTvxXF4XIDmCXvnAn1PXyxemwkTralf01YLFO3
KfekoBXt1lJAdIvRhcTAjlIIlXOKy52p0JfK03OT5IqdkQANO8sDMjiKqg6cEW2U
FnCbUCXaZnUD4usvP3W+rX3ZV8hsQBUktecC6Ic34HT0gaLbfNbKKZTRaSYN9rOz
mICxaMdyB8imW9lvN2PT3Wyeies9NHiEkhkRj8Y4i8cMnecKVCquZemh+P/MQyZy
0YzxYtWsI1G7lZPprym3FfftoxjPsicVjy5Wah0iNNwy1qnQc7nOFaKCGkp+xJjP
aDZn9736tpD0ks4jWgm4sHWSJSD9WgRyGdkoWYxG9OdWwL7IJ/8q6LqkJmJg2y2e
NN/VigZ0ygePbba6ET5D9H3f93QZeIU5LtgmJf4aeU2Wthm2jX7z0ifLFbtr8tuL
vCI3Bz7p0mSGh58bgEd6POFi/uD4Gh9B8/CtK9w3WbWr2ML1c+ryInREoEmUt2mZ
aFihkfbVwDQfukcOQpRjfmFzmPF2pSWhRWvrSkdoJ1aCF0P7VTS9JOOq7BJuktQp
pIsfQ8xeJcwYVxv37HXM7/q58RAnhujeSxD9TG5WRRlknGZfIrEMzo6sfry74gvz
ElgX/NTyx1DcHvZBO2NJVGEMJC8NnCI3acwJBJhJzANrrXKjUrw8nyXWfTDJTm7z
b55jggPJaeFG9JvIb8+NL7va8Lrz1baW+lNl9aUOqvNEyiubDRY6XOrrS/X7hICy
yw3JysQypwdrZuiAeGDHkGkAUXFNnwksd6lUEL62xOF2RYZurRMwcVUDrapBDarc
wH2JEUSwI45oOKHhX11XGWCdKvlx//VUof0Yc2bMXvLfJb164znreDZSbKSzAtFD
Rxnfrzn21uH8zMIYv/m3OsufpA5xrqJ/DZwoElEw3R720zcWZVccXWmbBeLAWpyt
I30oTF0eHdDNC1IzOPeGwfUJ3Xl/J4x7/raBBKoTQh6Qvd+5Ytyh8QP0NKffKGy4
u0WvdrSX+KmrL4lE29Bj59posp+BVl9cTb7Ex81Oc8ePc2Z5XU0lnqSY7y1vA89+
JpdZlU/DOnH02U4w7iqmET1QX1yEPf/U+m7l6mSkCUPd3EW9hcl0bdmChlE8k0lh
Yt1F2KPSwHR8vBO4FQgxIcwXZ1PlSyxMy7iDBzf2FNVtV/NsXtzXyrErVucQtiRj
aofMcUGwOSG99IWBy9QUVDMGmkUI+5KmXO4dHYMz011wgRiQATOfE7JLuJHJbZvC
CnK+wF3xLlh4N76ZtEKbfgIxFTPawo7a7Q1ZlZijVHlPVbpkkIVvbZ7/5jGy6XHg
07msDfBGsUz5dAfnUCvUDqPYLpZmUfZQLgS9Urjbiv068LS01hhm8+mOZrfwsdke
RMTyze7nfUvib6PhmviRKsjPdMAUDcZlaJZukSdv7c924vUIKojmtowOOsQs41p4
PQF6J7LWkZ4Jk/mGXUiM44Eds9GHfYW2hSqWc1fWS22CaK/pTnj7E0YV2IyZCJZy
nlaHhsV5GY4L05mPNcJ08ISE5It2hiYbO30INQi/gazQ9KkxMlEv8tjl34+3bENi
B+qkjgCSRiUinNMNIB+z9R22nptP7z8i4D7jYuju9po71ugbzCEPZjO6Ix/NxtCb
`protect END_PROTECTED
