`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MfPjULuBb40WAr9LbE9k/IjHmZxPV6SJYrA18CLMc86oHDRqZ/4p4/yNdhvd3FF2
yFYeNn0GVhSmtEdqQCG7swjpp1yUTqglXYIj2eF3xuruoSqe6L4nZARJSj9IFDvE
Nn4mDmoqpycQIlh3lxWcgyJMhLBaWpEg3mlHPl44y4ylmpm8S6V55YlOLYAN443l
k6uMbaUs5/WZB3iPJp6NOjY+jB7ckppwMFrZEUIXlg/m42tIjt2OK5q8pws6jtOj
m3nJv58txxyzno45VCS/F9QR4b1HO7lHK46+9hkewqJjqZoGF42zPuF2nLU2HQof
bddHS28SqgucgXYOc6wEBaN8+chy42uuAO+JRazs66Daz2ay4Hg63+iJXViA62mo
Wnc5qrrIl8EAJwu2Zj9Pr1ACjD4y38OclDdFuBwXGy0aUSSNMsivv99ZUpxrHK9l
7nz57D9BC8ltJ8Dy17IFaAt93gw/ixMAV0E4XERqsxltllBKzPbmhJyRp2YbMYuw
i7ELquBUohfyy+uPogXHDSwtpuWz7Hjt3jnh2fH9qwsMK72WFSR4Btl0anOKMNUH
ECAesczfZ4bK+bFDI6qSoqgRbJQ00tTxTeR3fnSSpriSxQ+ejVqzOqjaZ3s062cF
syAMn9G17jUlasu8XT0QQCGtp/R5NbEDYLmV1f098/KFer5tkP5rqD5h7swH9wgc
Gz3ZnHvMf21d0ynkdn2sPRtBkswlHmh+SdoKMbicaCLlRynUXT+L3yMqNfGWIzPj
9BQgSRzmVcPaIhaXTh/eGwE/TAq7zEDTQotgoc7/Dum+qxovGXfsunlCf8WTzjU9
kd+KpR70Oi3sqonV8V28cNFHT9+6X1kaaVpXLuDJWNlexxRoadi+iwKWmTmyzMqo
oCtdKwy87mjydA9VAkKLcGyru9pMtXAKOdjXUwmFXgrJgmEK8Mj8pU8EA9LO/VJ1
lRohUdwwFD2cOnaF7zUVCew2t1y3RXefPOWcyCG6pxUhTgys55ByMXqDlPSCszlx
iliD3ZrmS3uoYuiGBFYHbYK9bAzW8eMtqRDSG4UKOZ6b4CQTcq1nW4KFUP/yAYBt
GJxtI0R6IKnAOT2+jHqw9k+Pd2gSh0xO5ZSvxvwJgXICL767LnS/T8szBwrWL4BS
JwkXRGzAsrJJISayrQ1vAcEtGN5/4INIpNIKiZKgLzoYSPUf/THxYq+RKIfsMVG3
yRh4g28za4Gnn08SiMG/ncJaKVtN37wQ7cUYeR3CVnFdrYvHlOeXJ3yRYfuMSr4E
d2CbAO13ozPbebsxhRRH3WsahXaz1X+++DIJqtvR5WD5QjkM+FtLryH6/Vok6BZZ
xD4fDlK+Yww0hLzp71ZBkgO49kI4SzdBQuOyEEqrkApItc3Dybe0jFn6MDc7VCqs
M2hT745lKeom60gNUchVDDdjME+aBgVZPOqfahwxeegAZFF4iPSIKu/GkM8JLaey
DlhCxg2AieELPyL193aUidJHf7gl6Y/yUsnhywayIJpuX3JZzapBnk1qmB9hWinL
6JVZFQnmwT5S1XoYoVgXiRbzxydq4zyDrpcxMmcIYqPbrjO1GkiBO9Hh6pP8DNLU
fTfgI85S4Lf74iLVwumLftogdcvTh+IotPwimEA7gM80nGBllHQrAVOGgW/hXvaw
xVoT8H6C2PFq+EGEwaYFEjW7fSuLlFmfvzEmy8/IJjSDfrDeaHtHFx0EDSXgFmlP
H9KXausyGOZOs0E3aVlzWDixmkbGeyXd2/YUnvZjwPcKUx9Acsym52Uns0OtLtlu
mU44s3uovccslDaZU+9s/EEw13qDFqO1eN0r97swq6aA6eXx8NypFPiI0hXH+z0M
FFwF0Bd9Anhowc3sptkT2KrSz0jJ6/GVdTdzwif40+LutnH6mMxVLnZxE2fH0KbK
jufKzEFkyoyk7r9un4GtPKxetGSk+zg/7a5/d/Ss4OKiZWhdmZnwC5Nm/BC+0vJ8
mLFhsFRV4Ej2PNtJnxgYVhSURMVb95ZI/sromsS4b64xiqAJ2oSKgqVHM6FF0Mg3
4lY92PhDJTVMgK99FQ4yrDLpnIlSRzTiYNjLzFl6CVAlSX7mY+HrNJI1IWebrU6C
Cw3805M+E+oXdnVh1Rxoz3TKdODfXbFdvHlgpOgZtFlZZ9szbUweQO/tYfggNS/b
OaPL0HtEu9SdQMK221NAtNpP0fOtYEme8Tvtvn7k7P8tyW+A02HJWB4ydSyNB/8w
Du3uuxjQ5ooJNs6AYX8Wjj/1OW9nch2Y9JZdcU3BmmqrKREmiF/OpFec8WyHqYC1
HAhjfZBvfje+ZC8x0N46VZfeFDpSzg00PCgbbvLmbcu89Bza0qnZNMipeqJAJFmp
w1tyTtnck6Wbz+vVG9ucKG9HIxZiMy7HHX8QRuHe3zcoaW/6DaypDPD/BQBrpm1S
Soi7mubZmbtziuMawyOcLqmQxxxCBel6LwnXvZ88VdGniKUmhMuojkD1gITkfAo/
SPzy6+PPAaU4Z3t5dSNohmB6nmCUU2yndc/EkO6CPuv5s6uAQvL9OGsNBZUhnJDl
dO7NKSDUPbJMc0Cu99B/Kx08QkwmC+iTOk+Dy3KMyZ5kztq3qrljIlIhP6rLZSyW
YrcGD+lIHVGEV1l6bN/qXxnsqVZcGrP4hQgZG7mpVWAjLrk0vZx0gHmnDRD1pKsv
/VsOlQRFAWhaoYJkfD5qkz98DbA5GYbbVkBEksTtpq6OU8pzrW1co5eXnhkLBVNs
qvngttfZxWfEL0umX1D5MGmMUZU2KQSHXbJCPNjy+ez+u7mlslU8SbYAXgRHl2Xc
Fse03yJnvqxNnBN+lXyOXcw1+K3LykjIjYfuyPYB3SAiF8xABfaRGtOPcYe7shby
AURMlj7K6gs0S1hQLtSuZIJ4Mo8uicjdrhqMbbHrNEW38nHdIi2Z0nQ6nV8eGjGr
HUanx+/0lvcbo0u585gW1yBvow3Ppwqqw3pucojNiOBpD6O2C3zBzhOmqFU4aTRR
9kRWHsXJvTZazvB77+9rRIQXV7Ip5v4LH3WjryInNTmnddIL496jBPwPg+9EPmH5
3oiUqjPsxeenNaGXQcojr860knYclVjyQqdoQB0jXwZYm3y6RjCI76Gwbkds620P
vBWulFe6EPiIxthDNQV6WoNuH0yD1OPQmRtcdugnTnuqd4pGIKyXTZP3hu4B6jet
wpa2L70kew3q9gNa33wdTRHPLjm3pVB+AxTEP5ZX6pdNSg35xVDmeko8EIx8VOdR
DBqvPWjovkTafcRiCOwymazX3RNKjHNo5vlSEYpVaImxeLYkKmOfDYXb9Z1CtmYN
zODosxMOUTtpyzlcn9GCUTbpR8ysnvgek8vHiF6Vrc2wablNs/AqAngCAh2ZTuOq
PZEg+dDQbRO2791SgHHikGDyPmo6j57aHtdkF3eBzwTm2rO2hfPBe4NY4HVwr1LW
9V8pBkuBecHmqigOkKhRvZ2/bx/vKGMD+Ech3U/IxNO6KpD74D/60nmouA24bEbj
ckBZHw8eO4VdqW2v8H2NWXm/NU7nMEGPf5Iq1iQqcBGRLLcrh7wqNiD3FCmnT7Q8
vlQksRkEY9viN+ZRChvoqKprPUuSKzB/5JdgFMxXzXlnxy2eDhXboYDnWcdVpg6h
x1Y0kJ7Bha0lsL14hIOBqT0EofKNfYje9mWHOVJEJ92btLQUdc0iBpRdB/IyMdL+
ujo+VB1Up9mWB+0nDficAkUO2zd2TUaOCgxpdcGhOmatqIft3EtwAbFnmpxMoQ77
EwwAwwdM/JhZXZfbKKAr74IXQPA2m9XBQdpv6t7C81SvzSuT+IRcw/m7Pu4JqvAt
Sy88ZutERph78ticTiOQqdyBdA3FfOEZqlhJXs2KcsMO/gdrWsnIosgv6PiDT+RI
bRmpq4qJrdUOpcQdsXWP+IZjkRU+YcDWIx46WoPbN2iy4KoKYRx77D9lVKopH0cj
9lQIFc4t7s5+Bg01KO2JQhWQHomIqINWSIYXieSliIy19Q5xtjHncuzi9vt6czud
3iUMT1RjDuUZ6T1rz7MBh5CHOOpJc+kcby9R4+zs+xhWgsdzkdtC/IFJkUXkQqYt
8QuQWm+oQw6X3tgwDmwrAL87T6yVHY7qZXNIsEiv8MNmAq079+OXTRsikR2p/x4g
6FAazAuK4PStD02tQ49V8445o1cJawHYdc6uyCyRvlAm44E1Oxg/e2byzdBTB2Ls
ugw4vteZrYgdhtY2i3IzgSegpMJZfwlGA4lErDEoUtPZqyxWwU4y+MxxLwMNmw3s
TX0FDDRY/mZAVhSEAA8LLBzxtHk2EKcAzy0xbF/s7oFjkuKVSfU9FGyV+roDHkdP
8usVa+xxyyNsKp4Tm2EU7Zc5tvJHamZel9tnYBAHScpH8bGvOF2NKsqlbl1SPQZU
s4YfZJ2H15VfdGJvYrE/PnV1TL/0gLwMTw9INtggKYg8CQgQxi12SHYt5QfCBgUr
7LXmMz7KHrQ6B2zmrlNjO/s3Mwh46z/1hwBc+iszLva+rn/U5uo++Sm1D2209aRo
UP1WNyXeZj9I+51DXBHhsSh2rIgYcfQ4IVDJjBHYmVfPu23nEmexf1D7xqbi6K5j
4CvKxCQkg1Bmt9WJgyNbQikH6gXHQg1jCv/KY3h/KH8YJzD7R6m0z9QbXrmLawV+
DXJGvTMeaYO/JFmGDUXQkIWwTd8Bod+I00m0oNbaUM05mD0zMKDCYkhcyMHCd2fc
i12CvwCMyzBy7yzy8B1TgXsYHJ+JMU0fCDrZwVwGabQ4rrqq5wu0ohVewdg6a70X
qSanbBhZH2yo/CEozj0lswuzNUbYp+hwWc32UBNTN3iJfjKa5vYn8EBZBLULWguV
pI1ioNzyeqYRbDrRNi1wrbOUD6oxZtbhaEyoO/cnYMUU+l/8smc9ob5GLUti3oBM
VzXt8ohbqrzx4OmfLJdJZJ2dtMOSCsWlURhMMRThg5eiT7Y5eLPFlFZE0hx0HHPY
1X9kjW0h1csd+ac9HgJTSWiQv2F8PpkXMlN5PagXWvNzzya8TBHRzgpVDUxhsm9A
e3LGLIvAa+Q3XcI9VREikdxvPQXwvHs0hzcIZqEyel0dgjNkpyFUVw0eFCbS6T+4
6kJAHrrkYUAbprFXQPxZXfHfu5Rft1lpTEPVwKdZGU4c/dz3hdOvpOB+qOfZVtAE
FStKBwSypSU1hIe1UUblKptJAXHo8Lt1ruFDLmnakaMXIeC2AnwoCr6omScjEB+R
XpbWh399oFRIr0XkXlb+K0sb9rh582dfSagqmtdUlYu0MKXzeZNeTMNQ2F831u+w
U38UJuIMn+36bAgUzWRpRmZGKTNgnKXV53Imo5jPd918lKq/rQ5mg4udvTS01Z7g
NCHSlG2+9F2zdyN7FaV7+XJkqZE/jjjDeiCvhgPYZQ7UGp+DkGP3Na6488ia2n78
s1AOoSrv2abkUpfErmPwalYWmiu6AX4ddRkA4+LbLlUillUrzK7R5+FuJnnHSLlE
GnH/nSLMrTrs9yen8GXKn5gS+t9kFPe2VaTbBkKx60wpsi1m3pf87IpcZg8DX+aM
f4NBAdH1jF9QfCFi56OVOC6iXX3eBymZGfuzSXrEhh1Uwl0Vf/iKa6bYl9tF2U3+
jASmXh67deSWGfJNj9rsOoZigxGEYzIQk41HXWNVhR+finp3CQO3gURAadV2ue9O
jnUPEOIYqCn4Oo3fpti9qUP52/KiZZVkWBHIL16VRgdV+sirQEObwwOs0/wsF00n
K9wTJMcgBOxLwmPV1gKaG6FfFNkPRk35ckuFR7dRk+CNyGsvbCaB4VDUZIWjHU2+
fOUgwQflj4VPzJL2yP5HVIiU7ge5rVa6Gv2YLdUaJBk6GDV7R8vbno1qjWwdbK7C
HgaVDh31YGIrMOJASxaoPc4KKx+iFk8TsLF9NKRMWlFNXGi8BTjEIMYILXJi2Huj
bQCCgZo1/hPsye8Q6b5m4+I1SO6ki/ODqaTvZgjGWh7nTrwSFOdSCdLSLy7NfeRE
gDG2z1UgBQlafdYAXdcZw2WogUXRBFIyr/J/ljhKkbEY7rJv6Mbh4Kg/KrBUyGVo
AW0B3jGU9MXBMPjHOHjqqECXOD+W0ANVgr85jZGOTyibVGD5jgebNLFsXgN305uP
RlJqgU31kIGF9lhgSg2+jaXyOs+pvhmEhFGfqk+mUEqFZqt+DckeLRtGymWBc24/
lb40rPZPM6o220INzM1lPekcDWw5oZR+B5JXQaaYEXYdGT9kPMcZUkSsKxhdhx2Y
qO7btcz/EzL2NFup8pp1q78B5l9dds18GF70vEe/ieWtuBv5tfcdSR32qwjH0yke
d06eY5TpkVBpdmh4yMm+CVFYRYp3LlJ4d+dd2OTypaLlcXSyeyZqMZNAPoI0TxSW
SaIrSKWk6k5TeEgb+M6T2uP6KihUvysl2JCaCno3mYzpWgu5QZOgUm4ryZicPhJl
cJ1lgLNlIClzHoqk+YKVrDZD9UlEBc112Ty48QrgTnEztsUELgIlnm/Qbl9RUAbh
TqbSLvQbDHQtjtgMIhw502f05IC6rp2IAOPDiOxV5zWy49wWq7awpuaRIMmex6ns
86kGDJVOI0buaJ49OFF5jJSEC6KsuLH157ycTkX04i9+/N8kmzWuMckAnsPpxk9E
pJfetyV0tzQPqnvA0hywNK2AEFOC9yvB50ZeQxk1418=
`protect END_PROTECTED
