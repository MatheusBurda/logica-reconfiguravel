-- HSys_tb.vhd

-- Generated using ACDS version 13.0sp1 232 at 2024.05.28.20:41:51

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity HSys_tb is
end entity HSys_tb;

architecture rtl of HSys_tb is
	component HSys is
		port (
			clk_clk       : in std_logic := 'X'; -- clk
			reset_reset_n : in std_logic := 'X'  -- reset_n
		);
	end component HSys;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal hsys_inst_clk_bfm_clk_clk       : std_logic; -- HSys_inst_clk_bfm:clk -> [HSys_inst:clk_clk, HSys_inst_reset_bfm:clk]
	signal hsys_inst_reset_bfm_reset_reset : std_logic; -- HSys_inst_reset_bfm:reset -> HSys_inst:reset_reset_n

begin

	hsys_inst : component HSys
		port map (
			clk_clk       => hsys_inst_clk_bfm_clk_clk,       --   clk.clk
			reset_reset_n => hsys_inst_reset_bfm_reset_reset  -- reset.reset_n
		);

	hsys_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 25000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => hsys_inst_clk_bfm_clk_clk  -- clk.clk
		);

	hsys_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => hsys_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => hsys_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of HSys_tb
