-- system_0_tb.vhd

-- Generated using ACDS version 13.0sp1 232 at 2021.05.24.00:04:43

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system_0_tb is
end entity system_0_tb;

architecture rtl of system_0_tb is
	component system_0 is
		port (
			clk_50                               : in    std_logic                     := 'X';             -- clk
			bidir_port_to_and_from_the_SD_DAT    : inout std_logic                     := 'X';             -- export
			zs_addr_from_the_sdram_0             : out   std_logic_vector(11 downto 0);                    -- addr
			zs_ba_from_the_sdram_0               : out   std_logic_vector(1 downto 0);                     -- ba
			zs_cas_n_from_the_sdram_0            : out   std_logic;                                        -- cas_n
			zs_cke_from_the_sdram_0              : out   std_logic;                                        -- cke
			zs_cs_n_from_the_sdram_0             : out   std_logic;                                        -- cs_n
			zs_dq_to_and_from_the_sdram_0        : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			zs_dqm_from_the_sdram_0              : out   std_logic_vector(1 downto 0);                     -- dqm
			zs_ras_n_from_the_sdram_0            : out   std_logic;                                        -- ras_n
			zs_we_n_from_the_sdram_0             : out   std_logic;                                        -- we_n
			tri_state_bridge_0_data              : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_0_data
			tri_state_bridge_0_readn             : out   std_logic_vector(0 downto 0);                     -- tri_state_bridge_0_readn
			write_n_to_the_cfi_flash_0           : out   std_logic_vector(0 downto 0);                     -- write_n_to_the_cfi_flash_0
			tri_state_bridge_0_address           : out   std_logic_vector(21 downto 0);                    -- tri_state_bridge_0_address
			select_n_to_the_cfi_flash_0          : out   std_logic_vector(0 downto 0);                     -- select_n_to_the_cfi_flash_0
			reset_n                              : in    std_logic                     := 'X';             -- reset_n
			bidir_port_to_and_from_the_SD_CMD    : inout std_logic                     := 'X';             -- export
			in_port_to_the_button_pio            : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			out_port_from_the_SD_CLK             : out   std_logic;                                        -- export
			in_port_to_the_switch_pio            : in    std_logic_vector(17 downto 0) := (others => 'X'); -- export
			LCD_RS_from_the_lcd_16207_0          : out   std_logic;                                        -- RS
			LCD_RW_from_the_lcd_16207_0          : out   std_logic;                                        -- RW
			LCD_data_to_and_from_the_lcd_16207_0 : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			LCD_E_from_the_lcd_16207_0           : out   std_logic;                                        -- E
			dm9000a_iOSC_50                      : in    std_logic                     := 'X';             -- iOSC_50
			dm9000a_ENET_DATA                    : inout std_logic_vector(15 downto 0) := (others => 'X'); -- ENET_DATA
			dm9000a_ENET_CMD                     : out   std_logic;                                        -- ENET_CMD
			dm9000a_ENET_RD_N                    : out   std_logic;                                        -- ENET_RD_N
			dm9000a_ENET_WR_N                    : out   std_logic;                                        -- ENET_WR_N
			dm9000a_ENET_CS_N                    : out   std_logic;                                        -- ENET_CS_N
			dm9000a_ENET_RST_N                   : out   std_logic;                                        -- ENET_RST_N
			dm9000a_ENET_CLK                     : out   std_logic;                                        -- ENET_CLK
			dm9000a_ENET_INT                     : in    std_logic                     := 'X';             -- ENET_INT
			seg7_display_oSEG0                   : out   std_logic_vector(6 downto 0);                     -- oSEG0
			seg7_display_oSEG1                   : out   std_logic_vector(6 downto 0);                     -- oSEG1
			seg7_display_oSEG2                   : out   std_logic_vector(6 downto 0);                     -- oSEG2
			seg7_display_oSEG3                   : out   std_logic_vector(6 downto 0);                     -- oSEG3
			seg7_display_oSEG4                   : out   std_logic_vector(6 downto 0);                     -- oSEG4
			seg7_display_oSEG5                   : out   std_logic_vector(6 downto 0);                     -- oSEG5
			seg7_display_oSEG6                   : out   std_logic_vector(6 downto 0);                     -- oSEG6
			seg7_display_oSEG7                   : out   std_logic_vector(6 downto 0);                     -- oSEG7
			sram_0_avalon_slave_0_export_DQ      : inout std_logic_vector(15 downto 0) := (others => 'X'); -- DQ
			sram_0_avalon_slave_0_export_ADDR    : out   std_logic_vector(17 downto 0);                    -- ADDR
			sram_0_avalon_slave_0_export_UB_N    : out   std_logic;                                        -- UB_N
			sram_0_avalon_slave_0_export_LB_N    : out   std_logic;                                        -- LB_N
			sram_0_avalon_slave_0_export_WE_N    : out   std_logic;                                        -- WE_N
			sram_0_avalon_slave_0_export_CE_N    : out   std_logic;                                        -- CE_N
			sram_0_avalon_slave_0_export_OE_N    : out   std_logic                                         -- OE_N
		);
	end component system_0;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_sdram_partner_module is
		port (
			clk      : in    std_logic                     := 'X';             -- clk
			zs_dq    : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			zs_addr  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- addr
			zs_ba    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- ba
			zs_cas_n : in    std_logic                     := 'X';             -- cas_n
			zs_cke   : in    std_logic                     := 'X';             -- cke
			zs_cs_n  : in    std_logic                     := 'X';             -- cs_n
			zs_dqm   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- dqm
			zs_ras_n : in    std_logic                     := 'X';             -- ras_n
			zs_we_n  : in    std_logic                     := 'X'              -- we_n
		);
	end component altera_sdram_partner_module;

	component altera_tristate_conduit_bridge_translator is
		port (
			in_tri_state_bridge_0_data     : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_0_data
			in_tri_state_bridge_0_readn    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tri_state_bridge_0_readn
			in_write_n_to_the_cfi_flash_0  : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_to_the_cfi_flash_0
			in_tri_state_bridge_0_address  : in    std_logic_vector(21 downto 0) := (others => 'X'); -- tri_state_bridge_0_address
			in_select_n_to_the_cfi_flash_0 : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- select_n_to_the_cfi_flash_0
			tri_state_bridge_0_data        : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_0_data
			tri_state_bridge_0_readn       : out   std_logic_vector(0 downto 0);                     -- tri_state_bridge_0_readn
			write_n_to_the_cfi_flash_0     : out   std_logic_vector(0 downto 0);                     -- write_n_to_the_cfi_flash_0
			tri_state_bridge_0_address     : out   std_logic_vector(21 downto 0);                    -- tri_state_bridge_0_address
			select_n_to_the_cfi_flash_0    : out   std_logic_vector(0 downto 0)                      -- select_n_to_the_cfi_flash_0
		);
	end component altera_tristate_conduit_bridge_translator;

	component altera_conduit_pin_divider is
		port (
			in_tri_state_bridge_0_address    : in    std_logic_vector(21 downto 0) := (others => 'X'); -- tri_state_bridge_0_address
			in_tri_state_bridge_0_readn      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tri_state_bridge_0_readn
			in_write_n_to_the_cfi_flash_0    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_to_the_cfi_flash_0
			in_tri_state_bridge_0_data       : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_0_data
			in_select_n_to_the_cfi_flash_0   : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- select_n_to_the_cfi_flash_0
			cfi_flash_0_tcm_address_out      : out   std_logic_vector(21 downto 0);                    -- tcm_address_out
			cfi_flash_0_tcm_read_n_out       : out   std_logic_vector(0 downto 0);                     -- tcm_read_n_out
			cfi_flash_0_tcm_write_n_out      : out   std_logic_vector(0 downto 0);                     -- tcm_write_n_out
			cfi_flash_0_tcm_data_out         : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tcm_data_out
			cfi_flash_0_tcm_chipselect_n_out : out   std_logic_vector(0 downto 0)                      -- tcm_chipselect_n_out
		);
	end component altera_conduit_pin_divider;

	component altera_external_memory_bfm_vhdl is
		generic (
			USE_CHIPSELECT           : integer := 1;
			USE_WRITE                : integer := 1;
			USE_READ                 : integer := 1;
			USE_OUTPUTENABLE         : integer := 1;
			USE_BEGINTRANSFER        : integer := 1;
			ACTIVE_LOW_BYTEENABLE    : integer := 0;
			ACTIVE_LOW_CHIPSELECT    : integer := 0;
			ACTIVE_LOW_WRITE         : integer := 0;
			ACTIVE_LOW_READ          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE  : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER : integer := 0;
			ACTIVE_LOW_RESET         : integer := 0;
			CDT_ADDRESS_W            : integer := 8;
			CDT_SYMBOL_W             : integer := 8;
			CDT_NUMSYMBOLS           : integer := 4;
			INIT_FILE                : string  := "altera_external_memory_bfm.hex";
			CDT_READ_LATENCY         : integer := 0;
			VHDL_ID                  : integer := 0
		);
		port (
			clk               : in    std_logic                     := 'X';             -- clk
			cdt_write         : in    std_logic                     := 'X';             -- tcm_write_n_out
			cdt_read          : in    std_logic                     := 'X';             -- tcm_read_n_out
			cdt_chipselect    : in    std_logic                     := 'X';             -- tcm_chipselect_n_out
			cdt_address       : in    std_logic_vector(21 downto 0) := (others => 'X'); -- tcm_address_out
			cdt_data_io       : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tcm_data_out
			cdt_outputenable  : in    std_logic                     := 'X';             -- tcm_outputenable_out
			cdt_begintransfer : in    std_logic                     := 'X';             -- tcm_begintransfer_out
			cdt_byteenable    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tcm_byteenable_out
			cdt_reset         : in    std_logic                     := 'X'              -- tcm_reset_out
		);
	end component altera_external_memory_bfm_vhdl;

	signal system_0_inst_clk_50_clk_in_bfm_clk_clk                                         : std_logic;                     -- system_0_inst_clk_50_clk_in_bfm:clk -> [cfi_flash_0_external_mem_bfm:clk, sdram_0_my_partner:clk, system_0_inst:clk_50, system_0_inst_merged_resets_in_reset_bfm:clk]
	signal system_0_inst_merged_resets_in_reset_bfm_reset_reset                            : std_logic;                     -- system_0_inst_merged_resets_in_reset_bfm:reset -> system_0_inst:reset_n
	signal system_0_inst_sdram_0_wire_cs_n                                                 : std_logic;                     -- system_0_inst:zs_cs_n_from_the_sdram_0 -> sdram_0_my_partner:zs_cs_n
	signal system_0_inst_sdram_0_wire_ba                                                   : std_logic_vector(1 downto 0);  -- system_0_inst:zs_ba_from_the_sdram_0 -> sdram_0_my_partner:zs_ba
	signal system_0_inst_sdram_0_wire_dqm                                                  : std_logic_vector(1 downto 0);  -- system_0_inst:zs_dqm_from_the_sdram_0 -> sdram_0_my_partner:zs_dqm
	signal system_0_inst_sdram_0_wire_cke                                                  : std_logic;                     -- system_0_inst:zs_cke_from_the_sdram_0 -> sdram_0_my_partner:zs_cke
	signal system_0_inst_sdram_0_wire_addr                                                 : std_logic_vector(11 downto 0); -- system_0_inst:zs_addr_from_the_sdram_0 -> sdram_0_my_partner:zs_addr
	signal system_0_inst_sdram_0_wire_we_n                                                 : std_logic;                     -- system_0_inst:zs_we_n_from_the_sdram_0 -> sdram_0_my_partner:zs_we_n
	signal system_0_inst_sdram_0_wire_ras_n                                                : std_logic;                     -- system_0_inst:zs_ras_n_from_the_sdram_0 -> sdram_0_my_partner:zs_ras_n
	signal system_0_inst_sdram_0_wire_cas_n                                                : std_logic;                     -- system_0_inst:zs_cas_n_from_the_sdram_0 -> sdram_0_my_partner:zs_cas_n
	signal sdram_0_my_partner_conduit_dq                                                   : std_logic_vector(15 downto 0); -- [] -> [sdram_0_my_partner:zs_dq, system_0_inst:zs_dq_to_and_from_the_sdram_0]
	signal system_0_inst_tri_state_bridge_0_bridge_0_out_write_n_to_the_cfi_flash_0        : std_logic_vector(0 downto 0);  -- system_0_inst:write_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0_tcb_translator:in_write_n_to_the_cfi_flash_0
	signal system_0_inst_tri_state_bridge_0_bridge_0_out_select_n_to_the_cfi_flash_0       : std_logic_vector(0 downto 0);  -- system_0_inst:select_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0_tcb_translator:in_select_n_to_the_cfi_flash_0
	signal system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_address        : std_logic_vector(21 downto 0); -- system_0_inst:tri_state_bridge_0_address -> tri_state_bridge_0_bridge_0_tcb_translator:in_tri_state_bridge_0_address
	signal system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_readn          : std_logic_vector(0 downto 0);  -- system_0_inst:tri_state_bridge_0_readn -> tri_state_bridge_0_bridge_0_tcb_translator:in_tri_state_bridge_0_readn
	signal system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_data           : std_logic_vector(7 downto 0);  -- [] -> [system_0_inst:tri_state_bridge_0_data, tri_state_bridge_0_bridge_0_tcb_translator:in_tri_state_bridge_0_data]
	signal tri_state_bridge_0_bridge_0_tcb_translator_out_write_n_to_the_cfi_flash_0       : std_logic_vector(0 downto 0);  -- tri_state_bridge_0_bridge_0_tcb_translator:write_n_to_the_cfi_flash_0 -> tri_state_bridge_0_pinSharer_0_pin_divider:in_write_n_to_the_cfi_flash_0
	signal tri_state_bridge_0_bridge_0_tcb_translator_out_select_n_to_the_cfi_flash_0      : std_logic_vector(0 downto 0);  -- tri_state_bridge_0_bridge_0_tcb_translator:select_n_to_the_cfi_flash_0 -> tri_state_bridge_0_pinSharer_0_pin_divider:in_select_n_to_the_cfi_flash_0
	signal tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_address       : std_logic_vector(21 downto 0); -- tri_state_bridge_0_bridge_0_tcb_translator:tri_state_bridge_0_address -> tri_state_bridge_0_pinSharer_0_pin_divider:in_tri_state_bridge_0_address
	signal tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_data          : std_logic_vector(7 downto 0);  -- [] -> [tri_state_bridge_0_bridge_0_tcb_translator:tri_state_bridge_0_data, tri_state_bridge_0_pinSharer_0_pin_divider:in_tri_state_bridge_0_data]
	signal tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_readn         : std_logic_vector(0 downto 0);  -- tri_state_bridge_0_bridge_0_tcb_translator:tri_state_bridge_0_readn -> tri_state_bridge_0_pinSharer_0_pin_divider:in_tri_state_bridge_0_readn
	signal tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_address_out      : std_logic_vector(21 downto 0); -- tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_address_out -> cfi_flash_0_external_mem_bfm:cdt_address
	signal tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_chipselect_n_out : std_logic_vector(0 downto 0);  -- tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_chipselect_n_out -> cfi_flash_0_external_mem_bfm:cdt_chipselect
	signal cfi_flash_0_external_mem_bfm_conduit_tcm_data_out                               : std_logic_vector(7 downto 0);  -- [] -> [cfi_flash_0_external_mem_bfm:cdt_data_io, tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_data_out]
	signal tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_write_n_out      : std_logic_vector(0 downto 0);  -- tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_write_n_out -> cfi_flash_0_external_mem_bfm:cdt_write
	signal tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_read_n_out       : std_logic_vector(0 downto 0);  -- tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_read_n_out -> cfi_flash_0_external_mem_bfm:cdt_read

begin

	system_0_inst : component system_0
		port map (
			clk_50                               => system_0_inst_clk_50_clk_in_bfm_clk_clk,                                   --                   clk_50_clk_in.clk
			bidir_port_to_and_from_the_SD_DAT    => open,                                                                      --      SD_DAT_external_connection.export
			zs_addr_from_the_sdram_0             => system_0_inst_sdram_0_wire_addr,                                           --                    sdram_0_wire.addr
			zs_ba_from_the_sdram_0               => system_0_inst_sdram_0_wire_ba,                                             --                                .ba
			zs_cas_n_from_the_sdram_0            => system_0_inst_sdram_0_wire_cas_n,                                          --                                .cas_n
			zs_cke_from_the_sdram_0              => system_0_inst_sdram_0_wire_cke,                                            --                                .cke
			zs_cs_n_from_the_sdram_0             => system_0_inst_sdram_0_wire_cs_n,                                           --                                .cs_n
			zs_dq_to_and_from_the_sdram_0        => sdram_0_my_partner_conduit_dq,                                             --                                .dq
			zs_dqm_from_the_sdram_0              => system_0_inst_sdram_0_wire_dqm,                                            --                                .dqm
			zs_ras_n_from_the_sdram_0            => system_0_inst_sdram_0_wire_ras_n,                                          --                                .ras_n
			zs_we_n_from_the_sdram_0             => system_0_inst_sdram_0_wire_we_n,                                           --                                .we_n
			tri_state_bridge_0_data              => system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_data,     -- tri_state_bridge_0_bridge_0_out.tri_state_bridge_0_data
			tri_state_bridge_0_readn             => system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_readn,    --                                .tri_state_bridge_0_readn
			write_n_to_the_cfi_flash_0           => system_0_inst_tri_state_bridge_0_bridge_0_out_write_n_to_the_cfi_flash_0,  --                                .write_n_to_the_cfi_flash_0
			tri_state_bridge_0_address           => system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_address,  --                                .tri_state_bridge_0_address
			select_n_to_the_cfi_flash_0          => system_0_inst_tri_state_bridge_0_bridge_0_out_select_n_to_the_cfi_flash_0, --                                .select_n_to_the_cfi_flash_0
			reset_n                              => system_0_inst_merged_resets_in_reset_bfm_reset_reset,                      --          merged_resets_in_reset.reset_n
			bidir_port_to_and_from_the_SD_CMD    => open,                                                                      --      SD_CMD_external_connection.export
			in_port_to_the_button_pio            => open,                                                                      --  button_pio_external_connection.export
			out_port_from_the_SD_CLK             => open,                                                                      --      SD_CLK_external_connection.export
			in_port_to_the_switch_pio            => open,                                                                      --  switch_pio_external_connection.export
			LCD_RS_from_the_lcd_16207_0          => open,                                                                      --            lcd_16207_0_external.RS
			LCD_RW_from_the_lcd_16207_0          => open,                                                                      --                                .RW
			LCD_data_to_and_from_the_lcd_16207_0 => open,                                                                      --                                .data
			LCD_E_from_the_lcd_16207_0           => open,                                                                      --                                .E
			dm9000a_iOSC_50                      => open,                                                                      --                         dm9000a.iOSC_50
			dm9000a_ENET_DATA                    => open,                                                                      --                                .ENET_DATA
			dm9000a_ENET_CMD                     => open,                                                                      --                                .ENET_CMD
			dm9000a_ENET_RD_N                    => open,                                                                      --                                .ENET_RD_N
			dm9000a_ENET_WR_N                    => open,                                                                      --                                .ENET_WR_N
			dm9000a_ENET_CS_N                    => open,                                                                      --                                .ENET_CS_N
			dm9000a_ENET_RST_N                   => open,                                                                      --                                .ENET_RST_N
			dm9000a_ENET_CLK                     => open,                                                                      --                                .ENET_CLK
			dm9000a_ENET_INT                     => open,                                                                      --                                .ENET_INT
			seg7_display_oSEG0                   => open,                                                                      --                    seg7_display.oSEG0
			seg7_display_oSEG1                   => open,                                                                      --                                .oSEG1
			seg7_display_oSEG2                   => open,                                                                      --                                .oSEG2
			seg7_display_oSEG3                   => open,                                                                      --                                .oSEG3
			seg7_display_oSEG4                   => open,                                                                      --                                .oSEG4
			seg7_display_oSEG5                   => open,                                                                      --                                .oSEG5
			seg7_display_oSEG6                   => open,                                                                      --                                .oSEG6
			seg7_display_oSEG7                   => open,                                                                      --                                .oSEG7
			sram_0_avalon_slave_0_export_DQ      => open,                                                                      --    sram_0_avalon_slave_0_export.DQ
			sram_0_avalon_slave_0_export_ADDR    => open,                                                                      --                                .ADDR
			sram_0_avalon_slave_0_export_UB_N    => open,                                                                      --                                .UB_N
			sram_0_avalon_slave_0_export_LB_N    => open,                                                                      --                                .LB_N
			sram_0_avalon_slave_0_export_WE_N    => open,                                                                      --                                .WE_N
			sram_0_avalon_slave_0_export_CE_N    => open,                                                                      --                                .CE_N
			sram_0_avalon_slave_0_export_OE_N    => open                                                                       --                                .OE_N
		);

	system_0_inst_clk_50_clk_in_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => system_0_inst_clk_50_clk_in_bfm_clk_clk  -- clk.clk
		);

	system_0_inst_merged_resets_in_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => system_0_inst_merged_resets_in_reset_bfm_reset_reset, -- reset.reset_n
			clk   => system_0_inst_clk_50_clk_in_bfm_clk_clk               --   clk.clk
		);

	sdram_0_my_partner : component altera_sdram_partner_module
		port map (
			clk      => system_0_inst_clk_50_clk_in_bfm_clk_clk, --     clk.clk
			zs_dq    => sdram_0_my_partner_conduit_dq,           -- conduit.dq
			zs_addr  => system_0_inst_sdram_0_wire_addr,         --        .addr
			zs_ba    => system_0_inst_sdram_0_wire_ba,           --        .ba
			zs_cas_n => system_0_inst_sdram_0_wire_cas_n,        --        .cas_n
			zs_cke   => system_0_inst_sdram_0_wire_cke,          --        .cke
			zs_cs_n  => system_0_inst_sdram_0_wire_cs_n,         --        .cs_n
			zs_dqm   => system_0_inst_sdram_0_wire_dqm,          --        .dqm
			zs_ras_n => system_0_inst_sdram_0_wire_ras_n,        --        .ras_n
			zs_we_n  => system_0_inst_sdram_0_wire_we_n          --        .we_n
		);

	tri_state_bridge_0_bridge_0_tcb_translator : component altera_tristate_conduit_bridge_translator
		port map (
			in_tri_state_bridge_0_data     => system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_data,      --  in.tri_state_bridge_0_data
			in_tri_state_bridge_0_readn    => system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_readn,     --    .tri_state_bridge_0_readn
			in_write_n_to_the_cfi_flash_0  => system_0_inst_tri_state_bridge_0_bridge_0_out_write_n_to_the_cfi_flash_0,   --    .write_n_to_the_cfi_flash_0
			in_tri_state_bridge_0_address  => system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_address,   --    .tri_state_bridge_0_address
			in_select_n_to_the_cfi_flash_0 => system_0_inst_tri_state_bridge_0_bridge_0_out_select_n_to_the_cfi_flash_0,  --    .select_n_to_the_cfi_flash_0
			tri_state_bridge_0_data        => tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_data,     -- out.tri_state_bridge_0_data
			tri_state_bridge_0_readn       => tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_readn,    --    .tri_state_bridge_0_readn
			write_n_to_the_cfi_flash_0     => tri_state_bridge_0_bridge_0_tcb_translator_out_write_n_to_the_cfi_flash_0,  --    .write_n_to_the_cfi_flash_0
			tri_state_bridge_0_address     => tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_address,  --    .tri_state_bridge_0_address
			select_n_to_the_cfi_flash_0    => tri_state_bridge_0_bridge_0_tcb_translator_out_select_n_to_the_cfi_flash_0  --    .select_n_to_the_cfi_flash_0
		);

	tri_state_bridge_0_pinsharer_0_pin_divider : component altera_conduit_pin_divider
		port map (
			in_tri_state_bridge_0_address    => tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_address,       --              in.tri_state_bridge_0_address
			in_tri_state_bridge_0_readn      => tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_readn,         --                .tri_state_bridge_0_readn
			in_write_n_to_the_cfi_flash_0    => tri_state_bridge_0_bridge_0_tcb_translator_out_write_n_to_the_cfi_flash_0,       --                .write_n_to_the_cfi_flash_0
			in_tri_state_bridge_0_data       => tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_data,          --                .tri_state_bridge_0_data
			in_select_n_to_the_cfi_flash_0   => tri_state_bridge_0_bridge_0_tcb_translator_out_select_n_to_the_cfi_flash_0,      --                .select_n_to_the_cfi_flash_0
			cfi_flash_0_tcm_address_out      => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_address_out,      -- cfi_flash_0_tcm.tcm_address_out
			cfi_flash_0_tcm_read_n_out       => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_read_n_out,       --                .tcm_read_n_out
			cfi_flash_0_tcm_write_n_out      => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_write_n_out,      --                .tcm_write_n_out
			cfi_flash_0_tcm_data_out         => cfi_flash_0_external_mem_bfm_conduit_tcm_data_out,                               --                .tcm_data_out
			cfi_flash_0_tcm_chipselect_n_out => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_chipselect_n_out  --                .tcm_chipselect_n_out
		);

	cfi_flash_0_external_mem_bfm : component altera_external_memory_bfm_vhdl
		generic map (
			USE_CHIPSELECT           => 1,
			USE_WRITE                => 1,
			USE_READ                 => 1,
			USE_OUTPUTENABLE         => 0,
			USE_BEGINTRANSFER        => 0,
			ACTIVE_LOW_BYTEENABLE    => 0,
			ACTIVE_LOW_CHIPSELECT    => 1,
			ACTIVE_LOW_WRITE         => 1,
			ACTIVE_LOW_READ          => 1,
			ACTIVE_LOW_OUTPUTENABLE  => 0,
			ACTIVE_LOW_BEGINTRANSFER => 0,
			ACTIVE_LOW_RESET         => 0,
			CDT_ADDRESS_W            => 22,
			CDT_SYMBOL_W             => 8,
			CDT_NUMSYMBOLS           => 1,
			INIT_FILE                => "altera_external_memory_bfm.hex",
			CDT_READ_LATENCY         => 0,
			VHDL_ID                  => 0
		)
		port map (
			clk               => system_0_inst_clk_50_clk_in_bfm_clk_clk,                                            --     clk.clk
			cdt_write         => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_write_n_out(0),      -- conduit.tcm_write_n_out
			cdt_read          => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_read_n_out(0),       --        .tcm_read_n_out
			cdt_chipselect    => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_chipselect_n_out(0), --        .tcm_chipselect_n_out
			cdt_address       => tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_address_out,         --        .tcm_address_out
			cdt_data_io       => cfi_flash_0_external_mem_bfm_conduit_tcm_data_out,                                  --        .tcm_data_out
			cdt_outputenable  => '0',                                                                                -- (terminated)
			cdt_begintransfer => '0',                                                                                -- (terminated)
			cdt_byteenable    => "1",                                                                                -- (terminated)
			cdt_reset         => '0'                                                                                 -- (terminated)
		);

end architecture rtl; -- of system_0_tb
