`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8JH5TxFhnLizhxtYr/yCshj3vit4egIxCVJSWKHsmiZ4rbOpSLwLN908zYZIX7zz
FGpvhJx79ssKGpA1DN6fXBervvmoOsCdyTUDLGlqyofrmClbaetZZQGcdukfrF+c
5b+eI5LBIQyBFsipZVZNyW0zGFRrZv4v0ktZhhHaAl9SMQ6s0sUjgAurTvzZ3Qgq
Wczo5dE5NwiBkdPE2OgcMvnJkYGqGxgxYKyeHZQvqkI720T2DcMUJ2ueFmCAiREK
UCcMFbgM9kJ6JorTEHT5WUr17ujG9VY23oO/mqiPgNxHCWQB7ujArmfDhKH9Jy8x
z+E/tGRDv3psNCZgthxUU1jpZImZE9PufSKFDZvwGyBrpgCMrLwqoL88NfPVCHR+
bqHKxUen9lq34QqlV70BOHfYERtJHXuBEruyuqarXUxDZU7ndlgtSNM55mM2VT4y
im8cp+trulAJ2XqL5ZzEW/Z/HfdPeaEe3uj/Zj76AbBn5eVS3m4zNAGwkzL5ECO2
8GovomzuLkOAN5H17XTxgNhiO2Y2ZPE5PYDLZy6fuR05Lfe+/4pH90jdWb5A0/3H
mcqPCb7c+3pFA2QRxGjoR5jeosAAyIk+jtVvr2AqfXIJ1aGjJ81whsZb4ejIi/xQ
C6rTUv8YG3Q5SasIgIbNrQFUi7VSeJLTt53qPQwWaQcByeqnIxD9tpxV3J7tqa4E
jtfsNYkH/ajNJ0Ui7IT9qGTtNvAtp8uFy8p5hz16UPILwKBfQUfrrd1UkXLid+00
C1P+Cm3StZGtbhoawmJn8h8aWugl5OPfjfXmGCsIEANYglbXf0+NQbAFA77lz55x
lQOHOp1kEH6n1umx/7CdA2Dr9qA6NScmBZGeWonCoZf8k7gkX8pW2LK4jt3G7BHw
msqx5L13J0jd5KABKFa6bPI33dZBqvN9kVbtbAOOHwGiPUqQONOLVaSdSma15cLG
znTX+wPPulSsQ/yPJUQs0B9dyGKvGdV976VXIoXZOSfpFYaGGYCcOggxfYb1PMF0
DzW7B0m2ymeqcAfSl6Xzn49OawJ4bXUAJrc4LVIz0CQAFBqJfNiRFgI8oK8gbaCR
PQvgxt7ro0N6rjgtLUJflIt4SP+anlAnlR1vSKYXgYVebp5Y9MEhi0saBNTS/f90
0tQP5HldjAeomMLaBQ0KJc4whjUyOIsOQhkrVKviMI/X9PRiRf61qvclT3eU2QnG
6/Y7qsXvXHjyLtEzfiiuoYZJsqXM05MgkwkVyBq+w14KHRi9MRLExs14kdbhMg1I
xtP2CyPYXP7g8xRa1dhHcivAvgFmacVRd9XMj3oqtahQJSrBEVaK97a+9NeFqg5x
bsIBlASu77gjATPYZ8qF0F0YuWXAdUhO28Ue6p36qElqDjecewJNQvFnO2Mgoe3M
U/HDE2SUWY7b/V1DSjcYKsBJEA1VW+Pag6TSpiqzXPV+IWXplx6EJCqiNiKpoxNw
MRnqGT3aPMv4rvqLWWjmu1/6TZHBL2IclRfs3Ge3MjhusEAAFHBoVU5pfgebgLrJ
9kBueAg0gJvw1ywMPkM0vUdpjfIhOVaKHZR/gFjZiHuqo+xxodETy2hPBKfO6HUI
Eo8biunVQrGuIiof6hfcc4YDAfq8mRMAA0hs+c+1ulReUNMRQ1pfUvCbEJkgX5fs
VsD34t/QVsZnOvucEnxAyVllO0Yh6Fj+x4MQnRmE65JQDcnE8jVdLSsOAwH0vV18
c7h88jbd4yHA6bjlh/w2JcA+IhNbZxXCXLFT6s2m3GwxqJu49/260GfePvyVYY1j
lR3vWi8vZHsK9PMK/oKB9oD+je0o2uAtJF6PEEs7sEjD05MB3JjUIVXrqo/8NuJ+
2kwL8Q38OFBZaVI5Ie1qUuozIOjyGhrBTVHt2oqw9z3wvrfQEbETavxyMybX5YdF
ApJa7t7QvtciTgbETJYPIEYeKZgsEWb5uWuZyoS64JIIseGGoSOwJoiGPL8C4lHg
lUHWh02xrpgsJtkfSKKAAoHE4eCzw2RLkbsysuG9CAS0y97DwovRNlqcsoVzcs3H
TO7c4gVzzxTPr/YxcY8tO/eJqX7w7hu4GIzluJtM6h1lAM5P1eETScfAcUaxjieI
mYTO/fIT02DCc6nTP/ifVPgtJw1Ioy5na4fOqH9iAY1uqX/ZLVfl9RGds9PC5Tf2
ZNWbzDM4Y8cLb7yfZhXIo7F/p356wZ63eJeZPOy8anwRspjDdZEIE3ezCeVSLYUY
5viLTECOP5KP5NLHqGB9JA==
`protect END_PROTECTED
