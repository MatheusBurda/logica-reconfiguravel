`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nvV/4tONgV4spbQ2yhHziBdcnEYHTthzd9WxDCXEayRVECyeRctG/dfCHnM+0VQc
PZ3iUmvTl3DMmqiOICOiVGDaEq7CF9wmwXBuhTXerDtfNZtc88ynoNla3yoaWoFS
K14nvAwBWZcWx8P7a64i9kKmpurzfZLaEcAZ3etAUO1ZLUr2ejLCsmqu039pvRDx
b8XSCaJm6kPszKil/Jk3Uo6ao75/5hKwNKyUjqjQQnQNuzdK+b1kdy5h8ZOXCj2d
khtKaAbRBOaNNTBSuTPN+xTO56UTMga/2F8qtOLxB0hU9YlF+PPnNdHDnqrEIztG
QQEZvwbNvE5BWUbCzwJ5yGXmFH7UTX3o/We4d1KNBN5Pvk1omdS1W1xeULggfTjl
jm7kKSMknF8Rh1ZUa8s44pU6u+RssmDEKACT3HOaUI+Ngurh+WF+tbULCqEHtfGG
EVt2B4AoIrhMAd+SjgY0x40GLB0mG6n7PsvxAamo2CTDms/EPSoWKPFEBgysZKRc
epDGQEcboL94LyphMY72eq2tB1YiWU2F4b5q8UcKiKZxDevDKxFVVivS8MdIOnVV
cfGEmE5JslppA4j/lfgq+L9X02fE7gg5wvUasDRC/5MPeTbfwCqXaDEZXx3fN9DI
YziByqovSDUE1kb2BgkRUASgFet+3hYww5esVddBiOOoBlmwED/+FA/j15jS3Swr
2KqA4O+vmS3SVIa10pghMBNNOShzeSWObAwyuDEd96M=
`protect END_PROTECTED
