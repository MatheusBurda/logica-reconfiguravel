`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TCz21OvGl4NhL4lcGc1XL3Jjo1Y56OnpmSBOvMu+vSw35QqnIpSNKrG5p1lC1UNW
4TNXXzW779Rgl2AZSq9FMJboJ65G0E0ClrIU5ABSTAcgq+66U8WZFsHZeMD1N2iC
Wp7g8b29VYQpJHe618wpN5aZ1azQKpaBWV9/xAgGFlBM+3A42k6OSFDENzbHWz/N
veGPDdYicYUTmdZmZ/zUw7Mu3pqEMsWwhnoRYpVovvh8D8i+ToJVcwG5Y4iApB7u
iHc2giEm+M3O4oFfmCS80P9uzpfwA/ux7Jkdkyb9Wgmh4irGpm4Gg2TpwxW9BUNQ
tg4sosWOYKo6vWFT4e7FisL7V2mx0/hOUz5F2eK8cr05X7ENASONUQKHJ6dkC5ua
YpbcAkU/fyyOdg/EdtPb/k/RiAmi4+hVbTCo5RsAQ4b4XiFtbC74i2TdLgryr5AC
X6ynmCAg+DmU11ICN8lltQ9IaCSVVNf/VYgInMud/GCncBf/NP+QCn9YifctWjA4
syxH+mZ2nvh9F1B6ZhNV7l5GXBqPe39wf/8y6gRaX3biBKFoM2J9+CrAnmufIdvo
1z/lAKs7bqR6ELsAANUseZHVP0bGKL30QpmMbWVMKuH6umXRLS1XW202jl8ySmj+
2/dScRKh3QI1QnqexZh7Y2H0YjNi+lf8aJovgeKTClCpf2HxLnwgnZyhsjWq3sON
61kSb0l5icTDOevtrmZKfmqrdgWOcAjXQFHP8c8XTp0k+N1r/sfD1F04ahlxaVNH
fv1QuR4QWaUowI1LMqZGbOowkqpzpWZZEz+Gt9bUU1ZlrujQiUxK49W9mSu8zFTr
Zulx7x6YYVuRWK599VmLmSFbH7TVauvNWC6PgfGNqwUP7TTJZttgVPdZ6Mi6cG5h
Ozp/pEM8L+xBW6eiVw7QsH+8rY9FI1LLEqtKOSH9fOIWMEHd7MUgQm3XSQeQFZq4
FNTMyfVSVvsYAi1NITK5zoXbO0W4Y3H2kPf901sC4SzLP7ug5fsxa8LjjdTSQj38
lNvTK+1nyhPAGBU2Sr26+jjFkTO8nodfqwDqqdq3t9ug1gZA7Rb8bXsYm4ChiazC
YxqujiT0v8/TMlw3KHtlSYxDyEBn6MvV/INaUr01mFAjV4RGFZ/gieDmrjVJ17As
qZ7IwjjHdxSKd7zwCJugkLuXrcxtxHRoY8SiD4Fw2e2ZTu147eOpk9KhaI6l+kqj
W39ohdZRfwZubL6YMxf2IfeNuTNrk8MIJb09ypDhWyF3qEQRb+Of2pWJZ1mmcdxu
sK8zKp5zgoh/DeJIfqwRfThJj39ee3kB7mkk2iY+fMDEw1uC7mRdEMIX1H0kyc+7
HRIAFwZDUsa+ZONFxXXx60YyQC1vigwGHbfkBy8qtbGIHc1ETR7EV6pGgRX7PrzJ
LDbMMDaKH+8Q09upL1oP0pM8x2FMuAQsCboq6ZpEfN82joLV5QrtQTQxvDW2QbGc
tVZbEITXWyp8lqqyFvcBJSuxx8xnW8LHZWDdeSEtY19G8mjhTr+tCvg7Bm6uQmvn
hXxmQd/Le4xAVae+2l+yBw45OceWGpCZABVwHHWGsy47KJfH4fymYkSjXTvcBjq0
qVpOCMBVQ3yPMYQCmS+u7iopDvGsPuCx1GTkZ0hIKKpEzPJT7V6xSoHIXWKzZiY+
9aAhvQUeH7VwF22B33J4WZ1r7t0A+doqpHCRYdLxeYueHVTtoV1MHene1dPQ3AFV
7TEfvoP5P4wfMOBsqK0oX1WflOafoRp+nf0ALQQQ59EnMvrfS6TLBq5t4UQ3IP02
SUIX7cxD5peHpc1GkYQ6WldOqlrR8gCw+6W3BicPejhAhtANTLj6+TtPoqKIzEi1
jX77V+J7vQaRpbBGU3pGi7IWdnss8PFoMvMaVuw8f32YzyXXFYk0KJo6TPIc7tdU
bVLDZMiewx4xihLEchi3d012XLoEreBvog0J90X7KBeBSTBM5kyX123dpTyEiRiM
XkQP0z1WhybQAxLd2mMyy2vN2v5e/J+1iwVuZhXcms1PuwbJHBQM4tGm+SXvtuCU
6vS7K6APWM9CCxg+C3g+c+jqoIUGDvBJqGZzn2fwKCNdpITdBaizvffk3IWta9l9
1b2iPkyWPQxIAlUicxQ3K8j6UmcmNMzZXqtKQnBhK55zMGgUU3ESVSAGckarNcHG
v3NpiLL41tIbXMcMsHGLqpNS8urEABjjtCcFsIUxo65IinibIb+hmw40aAxiMu0P
6P2B2gnRmU8Ji/z763uNC3dGWovCsKSGrHZubP7xLf8goQtCVWI1jOy/Ojcv0CSP
McQvnf2UfnUXVawz8cSAYtk/2weGmFfXym+8HctencvlAPLIAAom/H0Fpa3F7AQk
Ofnu04TwyDD/iw4dw8DItBn2h13mH09271PqzfrSvm2dD2KYxLzgP3bjNDRh475+
mlzkRBH6Tdg3URju1gKNB3FcruTP/tTwWR6PcNEfnkqv7XY8+YQLQBwpXH3DzAkd
1h/YUDB02ZePbrPPs+4//NcIEahX8VMGnere76JLoUxuZpU2SDSfprbBdhaHlvN9
vewCdu6sBkw8npF8lw0DfxVU5l5W/VEYX3+KaOOlU1+uEZK1aUG6YKEDinonsRTu
dbPm9oYyog7srMTRw3MozlSO5oBv+OZdwsc6NywSl85M2JOL5fFMmjM/nCErgmuH
9sQ0W7d+8WAqHt7agnYfdYWCR1y+AJRxMQMEEk3cHb32y38XTLH1TX5/2UXyyJEX
VKH1otklJ9U8G/MPbUVdbQURB4AxQSFiyTx4SzgxJl4BNoX5Z/BsA3BckgiFTOB6
bE7fHg47SBK/nb250hImeQ/TUV1hv3moxqODAbfdebNs8pudUw7xcrz3LgC+Kgyj
FtcXrdof2zNQhbZ3TH2XW3OY4aJw05xhXuRi/vaaDmaxZuENYztGmhoCElqF1qX3
fysLWKf6PGg+QLSWwZ1+Z72jL9kKSlwyKPs1++831P+nQZttlmE49cZ7x71FGFHq
SYfvjHlG+AIKpLWHhZoTDA/oMG4KT6i9Cr9XrVnsqGjWPUUTiPwIRXUUdQI3Sxae
YLe0YiZjp6qquwZ6El4kxoHneaBmQ7K2hcJViM6/YmY4SqtUrp9C7218MJkX0Phz
XwzR4VunQOBe95/4ONbne83tQr397fCPxQOZy3QlvvhSE4ER5XmCyBofS2LgDuV1
ccs5/FbrmyjGQcBvSHJjvN4nNECEvZc5kumusFYD6YH2CbI5psQa+JzQ+PunDh6F
m8HGI0cZQsXtfkYyxQZVA2oYdeokgL/ptvH5Ik/aZWpT6fnNvervs9rUaD6FTPUr
5+AgsBLCmXsYYlNvNKTin6ubMaqaLF0snvjyxEfJNPM5nIRCMd06tSxbqyi5Owc/
spZOcHdGBgcmH8/pxoY9iF36s4uiC30gyhozf63X1j0uEHFbiRW6+gaXBjlnfouP
eFA6P9nNUVA57CQwxpx1hc5Rkv/lvHfl2B+ilqur260O4etEUmdBrm0z1DRnp5HH
do6LNpg5CDthnO1BU6zksDAl+BxGfNE/k9Iao7g190T7AsOhbxpwavm25qUgjxYY
MmEBzUewtm9meN3xPwGqUIhe50BoYRDtisgfuM/2nyTdCMAjQgOaVQBTwh9sbDGN
f1e4pQwcC58bHAiUJmvROrgj0My/R/TcN04914GBRxE+iGk9l5Mwp/WiGVn72Zdw
wlCwrH2gj2+I1qUYqgA9omx1WdE+wNcLL7wB4bPRdNdxkymOimNkzyM5GokjmaX/
/2WZghjLlE93y/xbY4c4SF/fpX+5HJJ/14n8l8AnL2UOUJSI6dcV5+//xQuJUufD
U+AeIsdiIjRgU1x54PmCoZe0LSql4CpVVa/gQS1iLWAyeLI40E8ZS4Wz7oN/OM88
OwLNOX3xpukJ5QmS5mOCViFBBfwjs8qNCRKevwoncZ+R00C3wN9nbgBZaC0LpUXK
cCSXvfBoEo7WF3m2R0wU3OR/ZYLe2CvA5sHK6LJReUNj9XlSzZwgQo2sPAQhWpj2
MOQPevZQ7DjPujfrvJFq6zDtX17B5b3wJBGH+bzXOtykEmWQbPDBN6ODytjyIek3
nppJLU0NgNffVdptFjuZg5vFOuQQc/bOLck4xtX4F4KzsxjgzqTyXLMTN+ht4eZA
h7FhXcnPn890jjdRCgu70D/thbV+q2YTG8WBOyovSHrlLn9UjtToVnPItn4orKw4
Ywe1fzLVKOSDDE0sGYWhFDNu4kE2dxw6Zoar3bo94ayTKn4pfWuN8VxpOhxCnD9g
3YDJQfBx/CY8EXqCGeVgEd871r+u4JHJKfr6b+Go/V+Ur9SE948JjWzyHsT8aIDJ
a5TiOMILtVuT94T46kcPQvF9gCb+28NtVm94IjNF+IzqQZ8/XP2rZvCMY6oXEUZi
1ZdsS2nZDQSa0XBl/Rivd6ecR8txFtyCNI4HA46cD6krMSyFDDt3jda9xdEt+0Aj
43Y01NmeQPBsnC2KrZ0x3Sd6zvh4qyMuWLMO7UspkS53UCpf/TPSfVsBqYOreYds
33p3OucWvLTEBgqnkp5BAAthjmTvg4LyIzymrD4Xay5GKEzqEByXwxrcezWZ7h5a
lp2t6DAjG/72gvux5218XOQQ99n6+5Ii3R25uy8O3Ll9Ok7SSUUqs3ymFSd1EEn9
y9aFBFMwe9fNzTLEKqTN2cnHrxgJdPy1IttvUOENAPkYVpdhkC31l4UHC+STxu2s
VoqVEZA8LN/zXHdPbTSumGD/T0BgUEivSGdBgCCjYn/L7sBr+OAGPskuGtDAc7LS
uPOnP3Rm49R++JD5VBNd3df46FhQCKbcjljMLULo6ytY/Ipeu3ugnKNnSRy4qqg+
kb4c73H2MK3MiYje/M11o/KRhgedH8X/s6ETawEbmVkFPtCDvnltjkfOamTK9nK6
HIhzLtaC+Mfg1+HrzCLxkhGsBpjM6i8ECaSxsyBl+GULHNpbklnS8oyLRG2E4S6+
Wac3YnG/9JGK31fG2rHMqciotEPDgoF3A5Q5AOUQDtQjuZzw2HmQ07CO1PQH+LnV
wCsKxYAkZY1XfpFaBHLVAn0T3rdEmALuA4QTWldPBVjy12BaZWq9ZDGYTXsHO2ca
w6uySxIiqLRLsHgQ1H5MVmYpFnuQqTZjQZMK/aemmvvxWsb0/eO1Yr+x5msFZf11
tVNKbsfxDDO/2mUYBR2ZfaH+sjlaZeNRm/Innq+VWN+63EDluwsux02AzHVLvvvo
uceiejElSuf5TwW0nZ5WEnt/mu4XM4rHzKrh0P7E7ezWlLmbZy3bRcYAeCTVD7ai
DX2WFd/1Tsc/Gz5xLW7BFR0jvCqvIQzmWcRXkMQezxkt+m+jURzlzeYBRJq5mgEO
c67wFO/WzyqLop/QZqaLpfQ99JGxZGIsdQjyAMeEOYqGbtBTOXEBxajcFv2PHsoO
sUSUBNFM2xrgsHcUANynzdhIfyu0CluzqkQq5YlAFYBIzaQyPWcqBGY7Q/EJBKcn
BnOY4b/WTu+r7BnHljaA1zttu/zH9wqOp7SB2uJkYwivJlHjwGK3I6OCU/xapTeJ
/o5jZRH9f8SFx2wmIaSlsi/KXQhDx9wNsMvFpyqtfu92XQ+o71FAjnpnIgrOrMrV
6nGDEmPQahxV/w3sRFOyuSp8CkhWn6NoclUJb2X5ASctAko4H1fZ9N56mFWe+sz5
LAXYuWzJe7bFIx0JUqRtulnbPW9oSkKMjY5SBf9BCw+k1xZnCj9g9zTVQxqaFFCz
wUWqu99MxtI7LGMKIpn35Z2fkeX/dxZb/jD6KWk8ntmDZ+h1sscSTiZfsjxUq4Gb
OVyUOVu+Z01qhZp+duqEC9+TigxkeyjKfSa60WPFVKYr27QcrV2i36MCX4cBqSkm
I1Y/N7xVcLzwIQJbxs/z2xgHuPqK0wXMpBewYfXDUR2WxmmSJZQBqRB2x57B23CA
HE4iHkM5+WGRthnCFknaMs++ccHVaIzV7co+dWpr92GiZgQd4zJEo2mGzx15fIOe
UBW3YGsWRJ3xEggAbmR42vsJD/GJ3CBLDUCeclR+6/zSfggaTNqmuIkFvqnyhhVZ
9GO1WZpC7qTuOl1YHI+C0rOoSNLy8E5fUcvlTUTLB6BTQfPZj8r2zfiqPJpPzcFo
CpQnlD8XkpOSkf93CT1mMVU+UFr2V9A1L9RqQwHiDpqHj3LiyMpS23GUxEQjaqut
4sKOrlAL2g4vwln7hxNPN/WJMnEhriyNHc/ivqLdTViWKOHz2Y2vWiIjyKvQFpUs
CHHhejY45HigTZWrn7edZj5hrWgAKWq6H+ThOYggc4+q+BFtNWvt7FOotWn1MqPH
lvm4zLkNbotEZHqKrDoIlWaklYmYhf1kKaIEedNokV/xhgfdp2GkZ9Fc4pKyDZoV
XhZit7jlSR9295ul0c5UUYjkaD6LehgRsXxHjLB6CkCG93H7ixnKq00CotLdqZnm
E9+RyYTbUacTfqWVnFMNnM4SI/h5S9t2V2+6a4s5V3ILP1hmkjXhmp+bS4DL5dL5
ZVrBnui17Jio7g64dM40c4oD9mJ7nG2Dbty9XxLo0/FP/cZ0Kz8YMzGzkxQyNV+e
fZPR9COCF35p10oPW9DE4b+xXJDWF4q6Fl/SXs3vwtn8LbLMjZOFwdriH/vTnYOn
SlbArzxtqRfJ7u7K/6YUzWFhrKBS93iKzfSiNVWUtzxHYnRUekXIfybd+Rq2dHgp
lyAKR5jqtzuy9OIQKbcSZIAOXzYfsnQBo3a86LbpVRoMT0kUuG8RCYKJffrnba3d
m2BhPc+gGXwLafvQEpoFrIIHB+GOXxpmd1VEpQLkP5EnUtYnqLjGIBxcV8xi+xDB
GxN5GzH4wXLOwy0h+JijDVqW3bIhWaGajrEc7v493XqdNqECide1XlO4bfV+fSbX
p60pmcbqTLTR3nt/WafAeaYoAgkcPTFtYYo9vt8quRwn0OJCqtOiDjMiIxbks7od
9dzIoO3/00J83slSiLnjlP2sCquae9w24/2XZqLOH31goKzhlRNWQthDfu90MAOL
DbaAHvAnuFDcLdyscwNyjKyHV9hTSIJP3Rzgju1W1x+mX9c7lQ5nDv1fPHWC7FWW
Hjoj5RcH4MmoFJXY+V+gNVR0JzagssEanSdDiFPMqUPJ9hA5SZnvK6dyn3AOkIat
hNHT0EOd/nSscDVhwuV1XGyyMY7hkZki1YqGqa2J+/YhjDgZucHrlauW8JkyOYET
FxkMDc3rMQ6Wa2S1fDVtjz4yBl1fV8/ggxC52q2W8D0R2QnxxFdYq+hgIeZFIKmH
dglu49szqY7NYPQHsDxu82Lo04n1AjUV9GyhaAmQMKq3iH1rBhr4o/O1kCpCwLXL
KLmYxRyQa7zoQ2wSCUB/Ja+cyqlQu3VfFpSX9Mzxl51/JO2fjISjPeJ44sUztJdv
pegLUuUIG3/CPVu97WYmegn+SFHeVLQYHDkwTu6AoSaYODeLOJwdYKvk/TbKetJ+
TBIm6c/4WghS0S/YGYmoOH7x6yv5ZEMciNwSmNWZugr+px+3YnsLtqsPkulRlaax
AOLBIwyfqgj7cAIzRQPNccr1j/A2R6EyVanmjXsa3wXXqwedGpvLfQt2F3unGNGP
2EuP4g9QSNisPZDL+FG1YViEYYhFj337ne2NIeEHpIVbqnzla9GANEU7PJmglwXJ
8aYI86EWcw8McKWmB3m30DLBXbxxNEejPrN4/BTlpC/Fe0QchD9/1FBHTEBCBQWk
su/LUwMBHmY9Mq10vBKpiBQ8gdUW8anrj6x0rJOXQa44/scvSFhemD5oc6t2hJcx
yEL5hHs99t55ti7QltPhmZ8HV7NGZKWVHFL1duZe6ULZwHEF2CUpDPqALWXOsN2Z
OaXf+7kyAKM4YLl8FXhLWKbhekdU13CPH+lSnzIi0MMhUFatz/kVkpTd0PcK2VSa
YwxLQOrSv1jQvX/rB05sUQHGYAK/D8RBkDMgVNzOym6eMEsGsjPxAD7GTOgRxrZq
om5esCfHcAKQBQ8C7HOWU/+jzfFspd91XYjeqoq7trwGxCTTdaWa8KOM73AgQCPM
0sdtHlfKuHHQsrbWfdJBGtA9HMBjYbM/mfdp3P59b6cAm4dkY/u99ap32bnVssQK
NQkHqgyx/DUY+gL8cmfWpbuQXi0ZOQMhcgq5kh6rqM+mDQErIAaWUD3YwtRDR2Lz
FFbqVciHe6nqewaDx/xriUAeTzEcGPste7wL9wyze1AZIxv/FNKY955gIDX7LwT2
fdnmbIL397tz2Q14AIdowpNXErs4cdWlgFxgRaxLhJs3SygNrnnQJvjGW+L5raw9
OwS/Y1S43HHaQ8IKWZJDn5p/SNlQRH1lVg9A5aJLHFs1/LvH42xFNBvSRWxjZyxh
X1ehziPAAE0qDNMkxbJR7ocjui9X266C1IYJrBGbL76mX/UJtF5ZRoWRCU/nuMF8
vOlgE0qZSFVKp9FA4aUHzYnXdWGiKoRVp4Lr4vK2MArHCDuoCKt0tA1FvoIsfzZF
glh2o/IC5HJbpTz8vVrcR8yJLG2VnCDZRdk0/OfF8QU6q+DTDDJoO2H3NoB/MJFK
AtwIaNUthN9YKNhJcp9UTSGiOkQHj2iNGuTsNddidNRs/E1QP5W/nnFjaSt3UwH3
wuRzkfPFIWwdvrkC1GrzE1CW/Rj2ZA12I9c1rPXhLJQ1c+NadQa+fDReC6pjOryd
oSEEUKfp+RxCSn1Lq7mxcgNnN560uJGpXemK348GQ6ZUDI6s6MoIcqgNEw829c0M
rU9J2ygQ3Gup6S+tN08j5czcWC2ocSrtkOLCUfozqIm8iTTFqURUQzQkBA08E85L
6o8Q/4RJ4DGaOWwJE33fpLGp2hVguSOksZOlnETUMgr355x2G+5344w7JoB9D/Jd
ERpdg4bN3Gc1IvOSPo5cXsNDDDeWmFmC0k27XvRCSrY=
`protect END_PROTECTED
