`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rOq1zIIdypjghMSE+EPjMI9E1UbY69aOxaCjNbnTi1/msSmCZFTUHHiAg0lvSKPA
ScTncw8nttOXdIQ8AQF/k7tYaYHlzzyaGe2rEAXJxkcFQlRdigwgswGbU/0ZmSk9
UPOzb7kWcNq19l6i958rPzBCZYhemspjtqVNr7YQf83njTdCGxf5MlOrGYERBZ9n
PA1OhErU/n38rYmkoh4KqqnRZMeOueOMAfMTZTx7Q31VmcZSnFEkUU3BeZ4hXvbi
4GBzMowNpHpPinrJFGYAPE1aflLtaPgd03aux2zL8ZDv/YlQ51HH/suaMR9nx8cN
s9YgoOuW9YHjyCKhleSmmyHCnuRveLD/5QwFa5KjJtKvzKQMCJflcNYrjwBlWt8D
MnuNnU0P5/iOluUC4xxKdkg5S2mH6cvsNjFqnOzAQd4KtDs7ozM7iHK/1w4dmz+j
YamUrGwwnXfhpfzMiHGcozDGu37XY4hIEMWrJ4CXdhlWPQixsMmmP41uDgFL7iI7
ycfiTuf7VribtAFm7rfq5J9fuFRbDGFuEiJD+QYFJ91CdTaCfEAMuszD4KPBavh/
K0ZxDZD/kBEtJUNncKNS/COvr9BELg0D9iKZpMv6hONBCWgCY4e1Pek2k44ABFBC
Yq1je0n5tzodmYUZ3rvF18+eUnGIDV0q0bmeZnBD8I+UOCfiRWlHgtHB9L3mEtaS
Pwi9qQhTFCd2Dlq+bK/VxJfolMYogf7IvvDX5X/5wEDaC4VPIdMx7aOyrR72MQzZ
DKwvhsMA1Go7w6xOt/6CGYVBGYE1v9iwx1aibeWwfIUkxtMXyzMMvYrqLhF56Dlz
GSpkBCctRRYyuw8tfYC5fpUMvb0WkoOJM8kyCQ+fqDN+Ral7HRZUNMzIul2b2b3B
r9h9+J7etj/h/BudC97PMBOYyiRKi4ubel37z4s4Ec1Dyh9k6KjzU8HCpvUZsuRF
lKIjhG1Wh3lltKveaxvGcwn7XS+DKKaW9XoZcD9yY4IPaRhJ27+P8u4ehRxbTK1H
OkVhjRzeYsI2eU3+OuQBXPMkThUffMyBwEOm41xr5/10wLb5DCvAgiY6Nv5ZBBGD
SVebxiPiX83arQonBt9pac4x9QKZqAQ3D00V3QRAEJDXLIOdXP1DxyzEum/HKDG8
dTd68mAWROqn4B86wyyN51Uiz30q7+gmYOHco1Bsb39E6skEf7GeimfMsMO3qzlW
5tPTqletQ+4TwbB37c9uUvFa/hnpPyh0r6OZ8Uk0EGAAf/oa7Jv8S5iTSUVG2iVN
ivn3DqUBcNqlLtqfeuKa3bNaGQsiyOmWe8xY/zL/jg5hPWNC5Q8wc3YkyZLB9P8/
4nktbRz4N+2LOdUuWIxfNjVp/VidEu/GmREBPHZxMV6tskPlRzBeGOJZy3j/t6Ct
edUDG3W1wZ55r9XMBuRNY8P2JZ6Yuk2qxF5NGde8V4QuSKOjwW0dTK/3zQIjWiBO
HCMgayKd/+LGeJ6XBeh4mwi0sg4VnQdzFwaCNpJQHcE1bIjNchgcXRVX2a7oe22c
oi3BCpBhwYX7pu/HjagRmQjrkyz83Ab7U8Ft8ElBZHgjBqCEKuiAxTd3jDTt7S6t
Jc5Y3MhATIkcJThIQS5ziyhArKaUWvawT0UGLdvVTYLuIJCBs1cBd9dx8z50R6JA
TCZgyueZxU0yQCI0XPF2CLFeKmswlpVk6CzTc2bkLAftqKVwWmZxAz0vuGLzsqXO
PT423tRohFDytODKigPYg1yJKLg1U+UZPoGxygwXGCYyZwX3EBUVqml9bm8qyio6
QyPnv7OZXbzS3IqfNr8x7rXyx1sWMaXNQdSmZ2RQVMtSMAXaB5YRZb1PMxjdkUJo
2Xc1oTkK8TVtxqSX95BZfTrMU+C65m2ZMh6wYMbU8vvggbyKX2ksActFMKk1gu9N
ssTBGLwRCxFAf3YFz+LB6CXrgsoRN52wk3aBw9CIYVcTSy3VUShBlnPhb7j4ezWu
ie9B1Tn3YY90eP5pmh10q/XQRN8uD0c3ALR9bcheZnP+1vvcCTeWWKDCYR5pV+9L
i6tWwozS/yRLWMvdgaU2VEwNDLrimEE0dJW3oeI0Mv3LWcWclFf8duNodSKkHabW
A8SkiCw2EIXovm3Ez0h+oawOvcD2xamHGkrQa/OlbMxv1h5pXt4SxK3L9Ss8Bp2i
i9xCLhunlGCd3gKPkyFFU00FHiILY0T1P9sL+pSCRum819aLOchckEx6ptceaWM3
ZNgPBEUxDRtCdltuE4XX9JD1WflCgH0hQSiuTP4exvbpPzIMfx/W7zUPoRBHOCVD
te/UlVAo1M6bF8bIfZzO8ThPFN8Nei6HYi9zW1iRaL4y9kRXEKb4WVxzO2DO/0UG
UnNkFzFvilq773KerFxiZxksGZf5LS5ebzqR8Px5OAg+qlRuPdvZsswW8vr2chFh
hV4WKcUlv4Qxx0fZ0SdvpVYxNfAQeaLAVF/kgymI9s+pcDt1rwak57ieRiVsCc3F
v2EynI5NSokS/FsI26+otztxYmFpSnSmujHtXsgX3D+7u/ly4lxleL9Qj/+WPrWu
XJHRunCpJWvKrbbFb0AduzKuKVjqrT0uWKCstLnc0z80VBHlv374VfbTx57uPbCe
ziKVqzFaWCWPdgkjBTGRhLfVfjkFXk/7VA4v4Mr3dBvOyOt714YvCGXhmxywNjct
LqxNTzwS4woFktMbyLpnSA37SOpE3bLNjWN83/fcinZqvF2vy1WhbhA+6LTFGFEp
Bm5ggYP12CLRoKjoMwJoJKNyLCAf65kWnthNMbxyeNokaq5wNepTDR/4f5TIkX6k
G1PZFSPlSgJkD3zSDmjZbMjUesW8VRJJSDZct+CSJWRrokTH5Spr7xpUPlDKyMlY
3Owa/iq1jHLS27+C2Z9q2ZjptWA+0V7L739XWKzv2Djk0ELEolOpUywu0PKWuodS
UKcsKii03a63UXT+mVNEzWraWhX1nvG+K4VX+w4DqKmmYmFVa5jclt6Li1UU+PY5
p5HhaM98olBWnmaIn1lhK5Touqela1YBZkXoKIGHlu4SLWDlk7b6QYPUTMe/km6y
urKwuyHLWw+LbjgfAlZlB8uCvH2WW19+tVXMCOmcTVbDFbLp3VHOD6YSISSeJxjr
drvlaYA+oay9FRq7XbPsVf9gZbo5tR+GS4VLswjsBUPyFGkvHgMdFOr72EFGsNlX
U9bhI8vDOQiNXSnCXyBrTuPi2wKSgr53fnZ5y5BdyZr9BwYInLKKCul+CgRP/CHb
VZr6g3Thcvjb4nFcLlRu2TSq5TVWLho63ujLPNAit0ztuSVCvNyOZPC7nkSHE9Y0
7gg7acbr865UCNKcICs+vm8TJppphNY/quNKTXRTfTLo0LSW/gaREcYHBFvVPKyh
yjk7XM3i2Q7EkZSgIPtGFNJHqdXsUAbJuJ3evJEyQOm8ViUVHgqyIZKu9SVxtqmS
GYa5UXGsSF+/7tfblqavDRv9Rwpsso1hpfgYfzUwIw9XQR1pkTITFCIi5g2ceFY3
HujuEcUnJiIDid0g68Dix80+icaOns7RgJhJRHybKTOQ9FrDFcQUOl3iI/172ga8
HhArxib+w4jLR8Fk6M77v7C70SBvf4TTzTv+E7SeR3tbtmLrlDvz8vAhAH0H8YL2
1JiJpGFZHJv7wgfW/We/Ijm+LvLqftY36IK6PIkHWQv5/NQ0rxferSX3iZxGy2/W
yaUPepeiLYJiel8Q1yLytzvgfhZiGe1ZtgE/gxExe02EkxIPBzLmKGau3rF7cqrL
IhwhiZEHWN9qel+wKtHCMjquUg0Vkqivr439nRdvp4MO7vy2jZOoX9B+RRZRXz9i
N8T9sXH6z79XWD1/Gd7FgeKBL9EUWnAZPcVZOCm+6y9kHAZ9Age82iRSCYtobA9k
Ny/0HdULjuAzJh57dJCcoF2/K5cgQ1UGq1DWwwso6j0kDsefckbj6g+Y5MUudK0+
Ot2CYCxrdsOCsCirxF5DCw4SLo2AN0GnHwmW2ilzBEvhGR0LamnTD/GDWr3vd9kn
e1FI/eGtuyqJ7qDYrCLbNMB2vRQ5Mu7/rCFTY1ajA2na1OFkLsenuJy2B3Hjcd3r
2UHSRL/esuP6d6qaPoKES0H8wJj23C9Um4Mj98p5+6f5/7LAi+oA4X6OcHEHMrpp
ec60KiGzQPKiVJ4dD/v3yGdb/0rqMRKQ5Wa5b7sWU5LoX3UeHdh7qYO2b9zLlnyy
53mhj5iQSdMAHqjZl+fhZ3sBFQAs5V8V7P1bNzJI+ghu6vfprabFK0kLW+MwSPDH
pTggbNHSwBggMFXC4frKaAba5kXkrD6i2qOPYfZ2wACQLfAS5RNJ3q0nrMSRZBtA
34KOBwXZxMS123a3lbj3Y4OHi74IAf1SZkli/T6jZy6UVujHoLyByJVFLZSlYXze
q/bQTBZCsW+aQl5Q2nu72JV5oEFUCf1GtI8VIwTJNujgKw3KEf579A5F3pP3LITC
hbBdlgzGhD1XlZEuz+McImwZC7kAG40BQq3cYjjig1fi/aGV4xMiB67STL46iODC
OwBVQf9dUVaPHmaZFEyhasEhkj4o0OwdgrDYS/diSztH+mM5cVhMoNm5mKSWb76l
wErIvXc8KnCjzh1hecKTfqxly+TRY9nsSK1rTqIWPA+TKe31eSzWCCbkHVMLnsUQ
dEXg2kL1rlc/8/ECz5E7cwyMoN6Q2/mDfd2BuKGsgEjpKafeBQ//qfX5sDja1AFq
5WwOCW1K+dGLsJQscY658bVWNVSy6plXmXQdSouoWTOTv/r9nz+c9xSediHGv9ma
vfJu3bvqIF7q4klKBClqos9bwBRfeCgjCKSYRd4XsTqzlofhVzu75S3jJpDUGH9c
pszmBcd5ws9ZoADo96o7F8IA64PB0Mjjzzk8rzWUlyhqZFQpVwy77gMFYoChDrf+
1VvoJ+OZPmZjudvrHEbUhyBti+Q3G3dai9m9i6Qga71MNWtEBHY0iZTPVBqk6h3Z
wNnnhhewR+hySbNspKBN8EymCV3PPgKSBubVJB6DnRFrQnu11M74nKAL9j/GGmcI
2lFSu+WplflPLs3BUWPpVve7kTY+oCKbmgRzK2GWMUop+1Nlp+DtOxDI+Sphoxct
T5oTYURR7TQqosKjMW8egdTkvGnQebu9cHoUE+z45ZS7Pmfr4H5vUV+bu/twd1uv
qqv3XTzr28OLjo3cs0lDWW6/U0XmLUCQRxCeXgv9OnJOI8RRBiqAYp6SfFU5Z5Mr
dLnz3c8qLk8tFhukgEkkl/Pt6KmOizv9aoRu1/G6PSYr/YSTzUaagvbHLRAPwG5Q
tThigtDCS/tCg+Eu8ePCnoVmtySzeBV8p78P6nR0wZaK07Piaz9+wOlx8tzF+H7i
xbsyLdynplO3ulFLiLFBm4BGkct+Yd/rtBwyU86Aq3OVxYVhlmNsHnBnTNvlhLdL
vzU/136qXLS8wlEbR1CTFZJBk34PQLG01cfqr9H+9FsgM3mZajqGwd9mTePycKo/
IRgtSTGoRUMOPkbCvIUG5XVK+12QJyz+5AspM9uU0edWnM8qWZ6QG/4pYScSllcu
6sJc+GaV/igCnRQUwa8zpM/t6qsfliK54H3uxzUS9V2bt3zew7TBiRow6bb9UvZf
TA1W1OL6kc8HxatQMHh/lTheRzM/pu+l2DqwQ56vcMekCC6En9kTP0Bzx3aut6EC
bwuN6ijoOIZWmAyzhXVPOxm97KlJC31OZIF9SECPuXvpf45gS+zLXrVfs4rx+cqN
sr/cSUhlzRlNWSM/1ejSC2cqmV8AgEdXnT1eqFPIZ85X8uOs4jqq2IbqEK9OGHy/
fp/GWv+AIXzovR3Art/Guk50SG79yggM0+20hkkuGxfWM1OKPN5zIIFxJc9wS7Uz
LHE0in+Kc/qdsrbOncTszQVmkY1L+H9EIBVOunzEcrJAGYL/6i2jQO9QsIgNqwY4
4B8R9HlEo2zyXhpiRhIoUBRf8ptOtmEqZH+edC9U2g3AqZSQUvTd8hUMex+jDyT6
mubv1UmzFP4p1iL+NFBZPJPm3s4743BA2yfb2TCbP6kQWIAVzQt5TDSjmrRq/mHg
wP6rkXbELfVmQqrizIobeC90H3dOtRCqqCYJD86aeUWDggmn6xNnlEm88F8mHHhb
Za3q/hTu7oxnIQjYhvH5zhAIKSBvn0ccVRJLJD8YggaIEgbsj9hI3jlEESymS4vT
OZcHe1eEKD2HxymQ4nnsEL49R4ypDAE5JPrwo1rGaL5U96TRfJbCep6V/1VO4q6E
l4L3KG3DNoylLkUdKFRNOU6279WotYzjcJu7yclMht7rDvj/QJJLM2sjf+8LTZtK
Rngj3ZgDOSZvdi48awwQKtSPhHGTWoIPf9OKWH0joRcAALJIS7WLMEnZhIh7dMVX
M1qrN0ylhfMZYGrhhqX0CXr5YtpwVoPP9u3VivSR90I4aRtN7pf29HLuSLVPKtNh
USyBlx+TmKl/q/1j9lgEIgYCAoN+05R4xlozQecX8DlJaXq53FDxJJ6W26Y18TVk
L9PxsBukJua1heRghUAJEoTWmus5NPdjRJcnj52VpFmxwge5u0Kl+VeIewVKbscK
0HS31Fhel/AsFDs/8wUNozq0b+uHJrfyW1/f8N7ikxCom7Ys7Z97nJj2yvPnqRDC
oGdtN6AL/oAxu3/QqUm17x5hlGqeGJKUw0N2uaWrajjtwUUeVS0jHSursePq2TNw
cGrSH+x0uO+ktP8dPNNm0hn5syNSpcaBc3KUtU4XZs7s9NPhE3440WonBM2MwRFx
VBdtraRDbl7yJ92hh/4BdMSbfigDOC74D3gh2J7yTlmfFPWI/8Is/7YU3doCdUjF
enRx5bh6/NUXsZwXSHKg3CyKp05RELI7WSu3k4NWQHGJdEgPcc4SKWDYd9KH3Ewj
qK1oUuGizCE0KvlOfO0i5XBdm7TgiStGRTUxbwxyndtGWl3vzXkBEB7m83K2Y+Wx
qaJOf1speOht4SHE/+XQXLf03d1mkoxTkM9yvYcET/EFT0Ey91p/pQrD87pD3pP3
0tt9oKtrijgxalZPcL9yPU6wt8k69zLyYA8ZRUrMQKHDg3bwpXFirlWSGfsw0cKw
CmxouRA8Epv8K0nkc/tI8EBahcaZujtRG+QJGHRXT4rSyRB248LYFjlRx3rB5An0
IwCDHlFopik2uFY6wg5SUniOUlfNiXJ8n8RdUhRINdqbx2o7OdvWUq49mWppWEiY
sQAhNVBNiOibxZ2KvTs7zXihZUMco1MJQHFSSUG1uWlrvJM41PTTvKb+InX9lmYl
r6uLUkntQkQm8ffZuemHGeomDLtP0k5TlTRGEMMs8fOtaT9EY+PTdZb8zrBPecQF
xNIDsk1uvRGD7aqQJVxCwUzJrzb94S/KOBmKeO+7+FXYMOEtsWWmkN+k67xsDer3
u3Kx+qmwQFs1rLy8phrdInDyIn4w1NcTIWJJU49oMYrZQEkDqx3Zyu070vv2zqA8
qyyiTjoBEVF4Myph5xOODCIEQGAfKIGivMJLPnq8bBtkl3vFlAnev9+8+6faG0+C
jOFvU03eGco61xMwB8RbzU8SKXozqopc+1PyEtdX0wduxDY0vJd9RmKAQfbiX9Qk
9MfQTK1wut/nkIUP+GbEziwMkWeVcMofUtN1Tzw0ZWT4E+kwNs2gRjQjuls6+bzM
`protect END_PROTECTED
