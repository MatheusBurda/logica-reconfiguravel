--Legal Notice: (C)2021 Altera Corporation. All rights reserved.  Your
--use of Altera Corporation's design tools, logic functions and other
--software and tools, and its AMPP partner logic functions, and any
--output files any of the foregoing (including device programming or
--simulation files), and any associated documentation or information are
--expressly subject to the terms and conditions of the Altera Program
--License Subscription Agreement or other applicable license agreement,
--including, without limitation, that your use is for the sole purpose
--of programming logic devices manufactured by Altera and sold by Altera
--or its authorized distributors.  Please refer to the applicable
--agreement for further details.


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity system_0_lcd_16207_0 is 
        port (
              -- inputs:
                 signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal begintransfer : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;
                 signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- outputs:
                 signal LCD_E : OUT STD_LOGIC;
                 signal LCD_RS : OUT STD_LOGIC;
                 signal LCD_RW : OUT STD_LOGIC;
                 signal LCD_data : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity system_0_lcd_16207_0;


architecture europa of system_0_lcd_16207_0 is

begin

  LCD_RW <= address(0);
  LCD_RS <= address(1);
  LCD_E <= read OR write;
  LCD_data <= A_WE_StdLogicVector((std_logic'((address(0))) = '1'), A_REP(std_logic'('Z'), 8), writedata);
  readdata <= LCD_data;
  --control_slave, which is an e_avalon_slave

end europa;

