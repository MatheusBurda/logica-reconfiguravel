// system_0_tb.v

// Generated using ACDS version 13.0sp1 232 at 2021.05.21.21:53:28

`timescale 1 ps / 1 ps
module system_0_tb (
	);

	wire         system_0_inst_clk_50_clk_in_bfm_clk_clk;                                         // system_0_inst_clk_50_clk_in_bfm:clk -> [cfi_flash_0_external_mem_bfm:clk, sdram_0_my_partner:clk, system_0_inst:clk_50, system_0_inst_merged_resets_in_reset_bfm:clk]
	wire         system_0_inst_merged_resets_in_reset_bfm_reset_reset;                            // system_0_inst_merged_resets_in_reset_bfm:reset -> system_0_inst:reset_n
	wire         system_0_inst_sdram_0_wire_cs_n;                                                 // system_0_inst:zs_cs_n_from_the_sdram_0 -> sdram_0_my_partner:zs_cs_n
	wire   [1:0] system_0_inst_sdram_0_wire_ba;                                                   // system_0_inst:zs_ba_from_the_sdram_0 -> sdram_0_my_partner:zs_ba
	wire   [1:0] system_0_inst_sdram_0_wire_dqm;                                                  // system_0_inst:zs_dqm_from_the_sdram_0 -> sdram_0_my_partner:zs_dqm
	wire         system_0_inst_sdram_0_wire_cke;                                                  // system_0_inst:zs_cke_from_the_sdram_0 -> sdram_0_my_partner:zs_cke
	wire  [11:0] system_0_inst_sdram_0_wire_addr;                                                 // system_0_inst:zs_addr_from_the_sdram_0 -> sdram_0_my_partner:zs_addr
	wire         system_0_inst_sdram_0_wire_we_n;                                                 // system_0_inst:zs_we_n_from_the_sdram_0 -> sdram_0_my_partner:zs_we_n
	wire         system_0_inst_sdram_0_wire_ras_n;                                                // system_0_inst:zs_ras_n_from_the_sdram_0 -> sdram_0_my_partner:zs_ras_n
	wire         system_0_inst_sdram_0_wire_cas_n;                                                // system_0_inst:zs_cas_n_from_the_sdram_0 -> sdram_0_my_partner:zs_cas_n
	wire  [15:0] sdram_0_my_partner_conduit_dq;                                                   // [] -> [sdram_0_my_partner:zs_dq, system_0_inst:zs_dq_to_and_from_the_sdram_0]
	wire   [0:0] system_0_inst_tri_state_bridge_0_bridge_0_out_write_n_to_the_cfi_flash_0;        // system_0_inst:write_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0_tcb_translator:in_write_n_to_the_cfi_flash_0
	wire   [0:0] system_0_inst_tri_state_bridge_0_bridge_0_out_select_n_to_the_cfi_flash_0;       // system_0_inst:select_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0_tcb_translator:in_select_n_to_the_cfi_flash_0
	wire  [21:0] system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_address;        // system_0_inst:tri_state_bridge_0_address -> tri_state_bridge_0_bridge_0_tcb_translator:in_tri_state_bridge_0_address
	wire   [0:0] system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_readn;          // system_0_inst:tri_state_bridge_0_readn -> tri_state_bridge_0_bridge_0_tcb_translator:in_tri_state_bridge_0_readn
	wire   [7:0] system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_data;           // [] -> [system_0_inst:tri_state_bridge_0_data, tri_state_bridge_0_bridge_0_tcb_translator:in_tri_state_bridge_0_data]
	wire   [0:0] tri_state_bridge_0_bridge_0_tcb_translator_out_write_n_to_the_cfi_flash_0;       // tri_state_bridge_0_bridge_0_tcb_translator:write_n_to_the_cfi_flash_0 -> tri_state_bridge_0_pinSharer_0_pin_divider:in_write_n_to_the_cfi_flash_0
	wire   [0:0] tri_state_bridge_0_bridge_0_tcb_translator_out_select_n_to_the_cfi_flash_0;      // tri_state_bridge_0_bridge_0_tcb_translator:select_n_to_the_cfi_flash_0 -> tri_state_bridge_0_pinSharer_0_pin_divider:in_select_n_to_the_cfi_flash_0
	wire  [21:0] tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_address;       // tri_state_bridge_0_bridge_0_tcb_translator:tri_state_bridge_0_address -> tri_state_bridge_0_pinSharer_0_pin_divider:in_tri_state_bridge_0_address
	wire   [7:0] tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_data;          // [] -> [tri_state_bridge_0_bridge_0_tcb_translator:tri_state_bridge_0_data, tri_state_bridge_0_pinSharer_0_pin_divider:in_tri_state_bridge_0_data]
	wire   [0:0] tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_readn;         // tri_state_bridge_0_bridge_0_tcb_translator:tri_state_bridge_0_readn -> tri_state_bridge_0_pinSharer_0_pin_divider:in_tri_state_bridge_0_readn
	wire  [21:0] tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_address_out;      // tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_address_out -> cfi_flash_0_external_mem_bfm:cdt_address
	wire   [0:0] tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_chipselect_n_out; // tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_chipselect_n_out -> cfi_flash_0_external_mem_bfm:cdt_chipselect
	wire   [7:0] cfi_flash_0_external_mem_bfm_conduit_tcm_data_out;                               // [] -> [cfi_flash_0_external_mem_bfm:cdt_data_io, tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_data_out]
	wire   [0:0] tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_write_n_out;      // tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_write_n_out -> cfi_flash_0_external_mem_bfm:cdt_write
	wire   [0:0] tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_read_n_out;       // tri_state_bridge_0_pinSharer_0_pin_divider:cfi_flash_0_tcm_read_n_out -> cfi_flash_0_external_mem_bfm:cdt_read

	system_0 system_0_inst (
		.clk_50                               (system_0_inst_clk_50_clk_in_bfm_clk_clk),                                   //                   clk_50_clk_in.clk
		.bidir_port_to_and_from_the_SD_DAT    (),                                                                          //      SD_DAT_external_connection.export
		.out_port_from_the_led_red            (),                                                                          //     led_red_external_connection.export
		.zs_addr_from_the_sdram_0             (system_0_inst_sdram_0_wire_addr),                                           //                    sdram_0_wire.addr
		.zs_ba_from_the_sdram_0               (system_0_inst_sdram_0_wire_ba),                                             //                                .ba
		.zs_cas_n_from_the_sdram_0            (system_0_inst_sdram_0_wire_cas_n),                                          //                                .cas_n
		.zs_cke_from_the_sdram_0              (system_0_inst_sdram_0_wire_cke),                                            //                                .cke
		.zs_cs_n_from_the_sdram_0             (system_0_inst_sdram_0_wire_cs_n),                                           //                                .cs_n
		.zs_dq_to_and_from_the_sdram_0        (sdram_0_my_partner_conduit_dq),                                             //                                .dq
		.zs_dqm_from_the_sdram_0              (system_0_inst_sdram_0_wire_dqm),                                            //                                .dqm
		.zs_ras_n_from_the_sdram_0            (system_0_inst_sdram_0_wire_ras_n),                                          //                                .ras_n
		.zs_we_n_from_the_sdram_0             (system_0_inst_sdram_0_wire_we_n),                                           //                                .we_n
		.tri_state_bridge_0_data              (system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_data),     // tri_state_bridge_0_bridge_0_out.tri_state_bridge_0_data
		.tri_state_bridge_0_readn             (system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_readn),    //                                .tri_state_bridge_0_readn
		.write_n_to_the_cfi_flash_0           (system_0_inst_tri_state_bridge_0_bridge_0_out_write_n_to_the_cfi_flash_0),  //                                .write_n_to_the_cfi_flash_0
		.tri_state_bridge_0_address           (system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_address),  //                                .tri_state_bridge_0_address
		.select_n_to_the_cfi_flash_0          (system_0_inst_tri_state_bridge_0_bridge_0_out_select_n_to_the_cfi_flash_0), //                                .select_n_to_the_cfi_flash_0
		.reset_n                              (system_0_inst_merged_resets_in_reset_bfm_reset_reset),                      //          merged_resets_in_reset.reset_n
		.bidir_port_to_and_from_the_SD_CMD    (),                                                                          //      SD_CMD_external_connection.export
		.in_port_to_the_button_pio            (),                                                                          //  button_pio_external_connection.export
		.USB_DATA_to_and_from_the_ISP1362     (),                                                                          //             ISP1362_conduit_end.DATA
		.USB_ADDR_from_the_ISP1362            (),                                                                          //                                .ADDR
		.USB_RD_N_from_the_ISP1362            (),                                                                          //                                .RD_N
		.USB_WR_N_from_the_ISP1362            (),                                                                          //                                .WR_N
		.USB_CS_N_from_the_ISP1362            (),                                                                          //                                .CS_N
		.USB_RST_N_from_the_ISP1362           (),                                                                          //                                .RST_N
		.USB_INT0_to_the_ISP1362              (),                                                                          //                                .INT0
		.USB_INT1_to_the_ISP1362              (),                                                                          //                                .INT1
		.out_port_from_the_SD_CLK             (),                                                                          //      SD_CLK_external_connection.export
		.out_port_from_the_led_green          (),                                                                          //   led_green_external_connection.export
		.in_port_to_the_switch_pio            (),                                                                          //  switch_pio_external_connection.export
		.LCD_RS_from_the_lcd_16207_0          (),                                                                          //            lcd_16207_0_external.RS
		.LCD_RW_from_the_lcd_16207_0          (),                                                                          //                                .RW
		.LCD_data_to_and_from_the_lcd_16207_0 (),                                                                          //                                .data
		.LCD_E_from_the_lcd_16207_0           (),                                                                          //                                .E
		.rxd_to_the_uart_0                    (),                                                                          //      uart_0_external_connection.rxd
		.txd_from_the_uart_0                  (),                                                                          //                                .txd
		.audio_0_oAUD_DATA                    (),                                                                          //                         audio_0.oAUD_DATA
		.audio_0_oAUD_LRCK                    (),                                                                          //                                .oAUD_LRCK
		.audio_0_oAUD_BCK                     (),                                                                          //                                .oAUD_BCK
		.audio_0_oAUD_XCK                     (),                                                                          //                                .oAUD_XCK
		.audio_0_iCLK_18_4                    (),                                                                          //                                .iCLK_18_4
		.vga_0_VGA_R                          (),                                                                          //                           vga_0.VGA_R
		.vga_0_VGA_G                          (),                                                                          //                                .VGA_G
		.vga_0_VGA_B                          (),                                                                          //                                .VGA_B
		.vga_0_VGA_HS                         (),                                                                          //                                .VGA_HS
		.vga_0_VGA_VS                         (),                                                                          //                                .VGA_VS
		.vga_0_VGA_SYNC                       (),                                                                          //                                .VGA_SYNC
		.vga_0_VGA_BLANK                      (),                                                                          //                                .VGA_BLANK
		.vga_0_VGA_CLK                        (),                                                                          //                                .VGA_CLK
		.vga_0_iCLK_25                        (),                                                                          //                                .iCLK_25
		.dm9000a_iOSC_50                      (),                                                                          //                         dm9000a.iOSC_50
		.dm9000a_ENET_DATA                    (),                                                                          //                                .ENET_DATA
		.dm9000a_ENET_CMD                     (),                                                                          //                                .ENET_CMD
		.dm9000a_ENET_RD_N                    (),                                                                          //                                .ENET_RD_N
		.dm9000a_ENET_WR_N                    (),                                                                          //                                .ENET_WR_N
		.dm9000a_ENET_CS_N                    (),                                                                          //                                .ENET_CS_N
		.dm9000a_ENET_RST_N                   (),                                                                          //                                .ENET_RST_N
		.dm9000a_ENET_CLK                     (),                                                                          //                                .ENET_CLK
		.dm9000a_ENET_INT                     (),                                                                          //                                .ENET_INT
		.seg7_display_oSEG0                   (),                                                                          //                    seg7_display.oSEG0
		.seg7_display_oSEG1                   (),                                                                          //                                .oSEG1
		.seg7_display_oSEG2                   (),                                                                          //                                .oSEG2
		.seg7_display_oSEG3                   (),                                                                          //                                .oSEG3
		.seg7_display_oSEG4                   (),                                                                          //                                .oSEG4
		.seg7_display_oSEG5                   (),                                                                          //                                .oSEG5
		.seg7_display_oSEG6                   (),                                                                          //                                .oSEG6
		.seg7_display_oSEG7                   (),                                                                          //                                .oSEG7
		.sram_0_avalon_slave_0_export_DQ      (),                                                                          //    sram_0_avalon_slave_0_export.DQ
		.sram_0_avalon_slave_0_export_ADDR    (),                                                                          //                                .ADDR
		.sram_0_avalon_slave_0_export_UB_N    (),                                                                          //                                .UB_N
		.sram_0_avalon_slave_0_export_LB_N    (),                                                                          //                                .LB_N
		.sram_0_avalon_slave_0_export_WE_N    (),                                                                          //                                .WE_N
		.sram_0_avalon_slave_0_export_CE_N    (),                                                                          //                                .CE_N
		.sram_0_avalon_slave_0_export_OE_N    ()                                                                           //                                .OE_N
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) system_0_inst_clk_50_clk_in_bfm (
		.clk (system_0_inst_clk_50_clk_in_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) system_0_inst_merged_resets_in_reset_bfm (
		.reset (system_0_inst_merged_resets_in_reset_bfm_reset_reset), // reset.reset_n
		.clk   (system_0_inst_clk_50_clk_in_bfm_clk_clk)               //   clk.clk
	);

	altera_sdram_partner_module sdram_0_my_partner (
		.clk      (system_0_inst_clk_50_clk_in_bfm_clk_clk), //     clk.clk
		.zs_dq    (sdram_0_my_partner_conduit_dq),           // conduit.dq
		.zs_addr  (system_0_inst_sdram_0_wire_addr),         //        .addr
		.zs_ba    (system_0_inst_sdram_0_wire_ba),           //        .ba
		.zs_cas_n (system_0_inst_sdram_0_wire_cas_n),        //        .cas_n
		.zs_cke   (system_0_inst_sdram_0_wire_cke),          //        .cke
		.zs_cs_n  (system_0_inst_sdram_0_wire_cs_n),         //        .cs_n
		.zs_dqm   (system_0_inst_sdram_0_wire_dqm),          //        .dqm
		.zs_ras_n (system_0_inst_sdram_0_wire_ras_n),        //        .ras_n
		.zs_we_n  (system_0_inst_sdram_0_wire_we_n)          //        .we_n
	);

	altera_tristate_conduit_bridge_translator tri_state_bridge_0_bridge_0_tcb_translator (
		.in_tri_state_bridge_0_data     (system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_data),      //  in.tri_state_bridge_0_data
		.in_tri_state_bridge_0_readn    (system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_readn),     //    .tri_state_bridge_0_readn
		.in_write_n_to_the_cfi_flash_0  (system_0_inst_tri_state_bridge_0_bridge_0_out_write_n_to_the_cfi_flash_0),   //    .write_n_to_the_cfi_flash_0
		.in_tri_state_bridge_0_address  (system_0_inst_tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_address),   //    .tri_state_bridge_0_address
		.in_select_n_to_the_cfi_flash_0 (system_0_inst_tri_state_bridge_0_bridge_0_out_select_n_to_the_cfi_flash_0),  //    .select_n_to_the_cfi_flash_0
		.tri_state_bridge_0_data        (tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_data),     // out.tri_state_bridge_0_data
		.tri_state_bridge_0_readn       (tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_readn),    //    .tri_state_bridge_0_readn
		.write_n_to_the_cfi_flash_0     (tri_state_bridge_0_bridge_0_tcb_translator_out_write_n_to_the_cfi_flash_0),  //    .write_n_to_the_cfi_flash_0
		.tri_state_bridge_0_address     (tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_address),  //    .tri_state_bridge_0_address
		.select_n_to_the_cfi_flash_0    (tri_state_bridge_0_bridge_0_tcb_translator_out_select_n_to_the_cfi_flash_0)  //    .select_n_to_the_cfi_flash_0
	);

	altera_conduit_pin_divider tri_state_bridge_0_pinsharer_0_pin_divider (
		.in_tri_state_bridge_0_address    (tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_address),       //              in.tri_state_bridge_0_address
		.in_tri_state_bridge_0_readn      (tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_readn),         //                .tri_state_bridge_0_readn
		.in_write_n_to_the_cfi_flash_0    (tri_state_bridge_0_bridge_0_tcb_translator_out_write_n_to_the_cfi_flash_0),       //                .write_n_to_the_cfi_flash_0
		.in_tri_state_bridge_0_data       (tri_state_bridge_0_bridge_0_tcb_translator_out_tri_state_bridge_0_data),          //                .tri_state_bridge_0_data
		.in_select_n_to_the_cfi_flash_0   (tri_state_bridge_0_bridge_0_tcb_translator_out_select_n_to_the_cfi_flash_0),      //                .select_n_to_the_cfi_flash_0
		.cfi_flash_0_tcm_address_out      (tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_address_out),      // cfi_flash_0_tcm.tcm_address_out
		.cfi_flash_0_tcm_read_n_out       (tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_read_n_out),       //                .tcm_read_n_out
		.cfi_flash_0_tcm_write_n_out      (tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_write_n_out),      //                .tcm_write_n_out
		.cfi_flash_0_tcm_data_out         (cfi_flash_0_external_mem_bfm_conduit_tcm_data_out),                               //                .tcm_data_out
		.cfi_flash_0_tcm_chipselect_n_out (tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_chipselect_n_out)  //                .tcm_chipselect_n_out
	);

	altera_external_memory_bfm #(
		.USE_CHIPSELECT           (1),
		.USE_WRITE                (1),
		.USE_READ                 (1),
		.USE_OUTPUTENABLE         (0),
		.USE_BEGINTRANSFER        (0),
		.ACTIVE_LOW_BYTEENABLE    (0),
		.ACTIVE_LOW_CHIPSELECT    (1),
		.ACTIVE_LOW_WRITE         (1),
		.ACTIVE_LOW_READ          (1),
		.ACTIVE_LOW_OUTPUTENABLE  (0),
		.ACTIVE_LOW_BEGINTRANSFER (0),
		.ACTIVE_LOW_RESET         (0),
		.CDT_ADDRESS_W            (22),
		.CDT_SYMBOL_W             (8),
		.CDT_NUMSYMBOLS           (1),
		.INIT_FILE                ("altera_external_memory_bfm.hex"),
		.CDT_READ_LATENCY         (0),
		.VHDL_ID                  (0)
	) cfi_flash_0_external_mem_bfm (
		.clk               (system_0_inst_clk_50_clk_in_bfm_clk_clk),                                         //     clk.clk
		.cdt_write         (tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_write_n_out),      // conduit.tcm_write_n_out
		.cdt_read          (tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_read_n_out),       //        .tcm_read_n_out
		.cdt_chipselect    (tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_chipselect_n_out), //        .tcm_chipselect_n_out
		.cdt_address       (tri_state_bridge_0_pinsharer_0_pin_divider_cfi_flash_0_tcm_tcm_address_out),      //        .tcm_address_out
		.cdt_data_io       (cfi_flash_0_external_mem_bfm_conduit_tcm_data_out),                               //        .tcm_data_out
		.cdt_outputenable  (1'b0),                                                                            // (terminated)
		.cdt_begintransfer (1'b0),                                                                            // (terminated)
		.cdt_byteenable    (1'b1),                                                                            // (terminated)
		.cdt_reset         (1'b0)                                                                             // (terminated)
	);

endmodule
