`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gD98ufLGNWTZ4biNhS4vMI27olLf24yqxl8yC5rp5YgwJAF/UXmJzbMarn10FYJS
57/F5I5SBYaAAX/ystdv5TO+kp8jP48mT/DGc7dgZAqPeimWYYYF1XACktzvnCyF
u7Gg0fWBek/cerGJvv1jlPEj4DDfXZGsXUH4+mS5mNR8d1t4RaxCYLAP/udF+jaI
3xwbbuZ2Kcmwmkm84Bf0jLoqdvE7PeJTihUMCHUQXxzyajLb+o0qTb3h4kpaSzTp
aY+FdSxycWPqyzElZxfKwpOQEkdzrmZeVLeVs4cbFFQJe6C5Owx/Jl7kJDcG77tx
uHl7ymi1L+l/V8ttxlJ8AZ8B5XrXUDgyGK3AqeK/mBeHHfWyy5/xB8NZ6KmqqdcE
e1RaZRI9iHugh2gSXf/sYaV29Y1hNJF3fF4ZGh7KbezFlgdUHdJJ1ceGJkpEiGit
cekTuWvbC3fP8fkb3ddqs5W0XLa/9fBqhR4UmUAgZabG8N8pyxOVXTmxuIp6c7Jn
SYiuRKwVJyv2eAz4F2uYJWeRONkZJ+uyeh6Slq2w3MjWsyIMlfVA6PoxjB60Mi27
3mB7jHa/zNgIHqPCoH8+iP0lEHEKc0HmxbquRFwbZxxK9SvJItO9R1wLi2TKTNu4
EC6YczZFfoKtKtu+gw8X6KJUqP7pxKGBZ0aNEikTuOG5ks1ATvSeh9BHY02vHGkD
BKBGOdHJ5lj8nAY/GpqSNsFSu5+6E+xvqMNc5e8HRPJwxxA6aQRcHokvFisjLGO1
e82qjDT1+AePC+GB1vPmGScRkAZ5zyuAoGvd96rpzNWNnf9EsITu7/wTv15AacHn
2N+ky9k/aq9R8uvEbpHDuy3W2R1D1ARgX/HDMRLeJ3PeeN2RstQJLm2hoCsynLF1
JuHcYvbcdT6TWr1sKiEO2Plrdrhzi+boGPYWQuJkh39dSSc4srw0FKkqQ1SkUNXx
ahuC94OcqMlWYL+N7sdtIgGb0k6wrRGYgnfS0Lm75ur09qIGB9ste6VMBWtlxBZx
Agfasb8PsJWGjVSpzsKUSITaNtE1+7C0kTuRc1XBubbdfqZ+PpD+Dwm6mWdDaJWi
qUt9MWLC4ubq1zt68qwCEaIcq8xaiZv6lDosStEeTCi4uXteUsNazCj5L5ovr7sN
X9VafB6N0DI+AjLJHUz6VPzj193a4+eO1rEiFgLX+u40ylVCYQnk0YfxAB0Xentc
bm3Bdozjq+owu0Na28n+k/PTr3BvOHZ/8OV7V6pPhAHMs7v69z4iZY0kxo7tdNgi
JeEh9ypQ2FEuWX5Yyi6OEcTL5XK+1LfvsrRm4tUEFcMsZ5Jl9aIxHMNJ/GSYBGuM
QxPniqFtvFtlN9nR1z1CCdGmuL5BZTHD69uPwjdCQCBEsD3VedK65ItFC9l3KEon
rBwzhZaqbPDN+sdl2KO6DqaJNz6y7hJaohxwIxv3JYkAPNKTNOHy0yH9Gdp/5aHG
Nb7dRGOU3oniq9/C9P7GD+Xr3KRLqhr+I4izBIJMIdHhzLQ+XG8uVs40kJc8di8E
N5icsJQWQEFmni4Awm1ygt38f3GfG4KcE5SoutFKhR4HAOt4gk+dazZ+IuN9co3h
HhZ5gC7bS0ZWPUOdVk+UWjfCdnBtGNe9lj+KY/2O9xzxhiDVn48Mfsf3vQ2dKqm4
dCOdO+9xm6hMLRU+YpFfyzsoZVaSSk+GFwiwLI04ikzYiVdz92Odzmnz5/wnSRs9
ucIEOf3dJ15MmrqVifaPxfbYoC1UF7rNVKX7AZNsAat8P4kwGEiu17dpmjwvMQru
h793Zl8lfkX5+eMx4pYTOQ0irWkCpC3XtgX3oTlhpkFUNvU8W7vD6ifbhy/GU6y9
hXEbLNi0X6jhnVQX556SNifhRj2RmZlycHpxf7YJ3G8024YkErtIQES/vikSw2QQ
ni4DGmRKq/FmtIQFl78Ut60CivodyAFkRZDbk5wpKoA3DZMMDnGeTdaYCN9o+m9L
Xr0dto0MfoLU9mesTminrH8roKjOTwRS1aWhxyIkQ+2MPYWeodcBjgonxKVuJKfV
5K0Js4ig/8ijTRFIqG50ZUqsITEW2jvNbYq8KRaCHagdvvhcJEMeXaI6Fd8J62Gm
BksHJxpRx/8QUpSVWkXxVrd30PIG4GOkdV7NImUBIgyPVG3F7ICISIfyGPKgTWSg
iDCovIShUm1KjFtydmaVy0nfwUXLoDNAwT66wdkBfwSRqehfPLexEpX4xrnKS4Xu
Yh1j8dYEXQEV6S4NJ2PfjX/H+zwhU4QsjQjFRRdWtpOVrms6a9nrwwJYE0a4lXub
3cBBFy6b8vLWMvVKquax8UGNqYvgADYn944IYiC8SJkV0FHe5/8Vt0UJXLTGwiMj
jztigjFvoomA8vuINx5DLMAcQH8a384p/BCKQxBt4h1PcacL8FCC1HCKDbZb35t1
zYyav9Uy9YG9TBnvuXIO8N0UW11O5boRTODGxPoSZdpmU733Z8h1YmUQFKY+krxW
jDmbKqQMk90yCVclibarGsbbw6JZE8zQz3raKmEVBFEtrNcHcZU8HtYndRkLQr6p
wB2lpmuZ/xiUXvDwBF9zxjY9s1R0z4HI08QetDPOc0yC6WB9OhOiSg1s+o/vS19N
ps+kqjflqlQcgkDnKDCC5xW3ZjYwnXrIuZ84oO9EoIMHrJMDZFVpHrCfJqQNdX8B
7bcEmFuSqG/5DgNZ348JNkuod19cvYY4tqsf3U9fAunb2yeO0+KLCpgHW6Z1Uy7P
aIRk9n/9w20ZB5sNugcZiG+CQrQWaQvKycZGmpI+02JZzJX5vQplrzW3RdQVEXkF
ivd2/BjhcLMiEUDZt56XMv95o0xqUgFFyqa83thFBIGk9piez7HnZyztjWtc8vnl
1efaC6R0DgV8eE7ugxfJLzhjnLOolLdkUgO3ZMz4OjZBTNHO7X6hOdfjgCB1qFjd
kJBSvSROsvtE7zESmNsg+mwjD3f0Km92J+DluOM7k1+hHmjbolcwgcv2iLA7cXYu
CP2891+Q5ejVVmRuo4ehsakssihu5RGCKBU1PPByi4PIUhsrrpTj3WEZAptuVfKs
KSfN+K3KUs5ZRHa7Uv279OJNoaV4VE6Pf61v3pQ6n3cP96i4M3gTl2w9acdEGM8x
PlywcJv++xXbzNMXiRvyVUMlOFbVLDHW8OPLQUBpQnFmrs8XCgE7KKxlDEsb77EQ
Feh7iC1WXFP7u/9zHiJBXh6HkTpAZqKYB+OLySqd8qvT0gG0cB36qEJOJOsB6ufa
MVySiNyNthPvWplKZl66OVmUjLgSp71OrKIaLNW0GITQPGXYm3yf1S/E6xqPF4w/
iiiYaBcVj02407DRP4tDQKcfOFMjmNVx/eLKwOdXdGkOsmoIgUQ2q4hpJ3Bey7HU
X1gKrC7cAxYXA4OSgzmJUztGmfnfONtQU/HVnwYJ7kkHqpskvE6gidi6IaJ2TOTG
JXhJX5X7K+J8f9kL7b9k4BHh6gnqViIRrDyF6G5uiU4d2ukoQCfmNFDX2MiIVHOq
1rhF2omaar1c4gFrF402kSAVLe8yW1Ea7b/eVpMBUKvKEjmKyegsbnvuNdyiNnU4
IDRHnETKWGNKFiUSFXFB6MhEikngtUkguHAJb7A/Jnf6fZIDpUDl5w1+6u93M5AY
MEpFyVdSG3WfN0LggHwKqAers9VGjIDSYmsRjbcMZ6BSPd0kubiTKjUv50CpCLOI
a7F4WM7dEXcvOD8ZSc+NXzW/S4wxGDoKFnTYQ5yEbMZ3a7IyT/YyMw0slNjmIo/a
FVF29cuCtk1Vg6d/BNZRSn6BIAEdxygaLjnLl5EB/FT8jCiQyks4KKtD2RMdjW8z
mz8T1w9eQZAoSR3bphvJ7ZppRwAJEmeO6w6r63WRBobAJemXir9Fmp5xjzkTK4rB
gk3wOsXQwAcCwlLK9A/btKGy2ztswNHHz1wjox8pVHMoYt/xGaQxj1J3vA8I1IlJ
0uyszohiDoym6kz5Z2ayIbJBFrI5jn96Aq3zeoyxdgL96ad9zOr0vYCmzGyLX8nd
ljxmpZCEAEC4GPL0AgiV3OCfrKSaMNrlOu4z0AP42zQ2vqbsGfZHtVugrawAy891
PD/n8TKUMy8QILE1TEWoFF7WJKrQot9qZUcWqOKlgHOLIvRR5FKcLQBRX2VmkQla
PD5UBbGAYNL9pffXqd728+G0DXdCRRsjz50+zkEZQXJ9HOpXAGuRsmn1RREjxLIU
sCxmLUKb/vXUFeUvEY0chl+cP0JMDR7NAHoBNgSZTwht48rq2bT/sqiJ33Vx0ofR
NId3ZnLyYST3MDEWofxcJqTFkYU+bh87sjXV2wRjAg3XVXOULu/rdJD+7uAH+XDM
W62CNtgvgFly8YuBnmAsOlEqsGES9FF0f/X37BmNgmbyUYRoCEVFS5VysASnB7CF
XTTWsXYH+P1bFVjhrp6PEm8dJOm1NnXWPcn3C4vbbJWXRemh7BPGkoM8KUfDPApc
KmsAorLw6jMSurtyR6nQvJgVhcjHnB63DEKxpHgWf9AVQAPnRo7HOBWeYdRi+Ui4
62iZDk8fmUG16c6RtVAGUmuiDDa2e0rQXykR9vW/qjxBPziYtDf1PxaV5h92Rj7F
MmiQZczY6adoL84Y7xZrw+umrvF2Rz9BVkTksqoO7xVKJjEatyYEIWY6/YX2yPuu
r95ENHTGXShhCQ3xTZuEVj8dZfi55qpRJE3Q+N8xNub2TQMG5OeRVNcctgRFO3fN
3YcSaQTtBPmdE9KqupaPT7CXU+BNdSsSpxxgSeP6DpW4g7N/4bIJ/t3H3qp0lMPa
UyvHyYpwGqfPMJVkagPast1gV91yRN+KW/eYxO48GH2MBACtyEqdSt7sXdIgcu2v
VlU2U98zAJHft9qpLC/KlUkhuwQxOnbSZuiRWBrgT+7pc2U1onGpUMFEOzyZCzK0
cheXYHPbnCY36Rj6dq3qQfhgkimjRr0w2UyAWcPVRMrcxJQvSahv69AXpn4P6/Ye
teWKj5xZCf6Fz4q3kNRsKqTzCWaB83EfwtYTsfmMmxkM1n693iDBgQt7zkDUUA3y
zk7+X1g1JcbfOAIARCD4EebvtpNGK+b/9fL+JaAZleyfLBQyieZAvxVVkbFm75Uz
+MhFQkw4R9EAjWShzOCgIXsHxDjAHPpton+fu5XwM70etIeXMgLTvlHBrGCHeKuc
iJGEPBq6qqV1aCtQjEdB7REpzHEZiTqN+IYHieFP4j2RyB3Ymj+k10rQrwdHvcKd
nHQoAMhGpf56BlGUsxtDvy5+CwewKwFJ0VCv65NdlKpJpmXHAy/OuFjDhVd0RSVG
C3d5piETwjLjEMgGS8qfUsY07zfLhRjMrDW/XEd2NMZJSpPJ9RIjsNvjMHBjrer5
0RruPLoNXkwtSvap+2/nFdLFsqYvcfdzrcsQ+EtqjPGTMHig6IatKAtqo0PvZuXc
5hcGwtrVspRAPVmlQ5sK92sLAjjHwfqDhcw/qWcTsvlyabfO7W9U9VIdt1e9WG4j
ED1lBSzF2VaQMEA62LoTGzq7y7cuDe9Eif6aKWdyyA6ENR0yLaMHS+MgC6wFxjyC
8/XOlrRHi13AUKfU4BuCDhZMM1LScTAjm7JT8w9khmvLo2GKoBQBilRREGaDwOPS
OwaLP1WXt5E8lPV7scOA6lHRgqRE/pKyXgpNT9CL+VDSd68YTKxsuibwg6ytvLyR
G/d+wcTeugH7XOhzONqIi3s0tKiwWPUB+vz64W6SGxkmIa7tJ+3QPosVS62oM+CC
aK/HlBq2wSIs0NOSDmkv08ESSd+PY11Qmf7GwAxcCoPCtSlPn5A9VPtAkxZV/B2m
0NYTqXqWrLLGvU+G2uw6yMQ993CjlFsj2CAL3vlyUSXV1/BwP5m9E04hbDmN+lmp
Q2R/lqoW+dI5Jqv3F0+dXDVKsvK8LdBnLzN8CTeY5UZO3SWH1u4ymmh9Vq58rD0f
xAhLAA0IAidAceLyx9qkF07F009EJMjoT1kTVe1PSigNwSyugKQuTXeExf2PX7QI
CcMwN28tA0RgeDS+GMC/pMumjOh9gE3giEcbTVDMRt0=
`protect END_PROTECTED
