`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UAaMo62Y1Y3Mm6KudggRgwS4O+sWP8JH9O6yoHK10h4IGkI9g6SueoBN9YjmNBCe
NGObxssQtxGdXROtAU+m5VNT2ZKYkK41Exjk3p3h+htt36upz8DF13sEEw3VhBmB
uzbZWsZltXJQt+w9qgBIh3Q3WeYP1SIohx+D1I+Fis5udTp+5wqQoeVNFWQgLwO/
19DakUip4ZschrcIN+ry01wP9nH/GnqMy71kF98lf5JgJy8t05RVs+trfewiD2ZV
Cspfw9MsPs6j1TvQWyWgv4/bE13OmQHZNQuW2MePF4HVNZSohuSAxy4pOd7oqsPD
DTw7F45q7885uZdRKoRQfvWHYCIoJGOp6s0f3nnnXOuNAazX5QVlHWrQB7bn/DhD
WmtPAZgShSUIvLSyojEs0r80ctiCaTpqt3iO+k1IVszQnVfet7n15j0i5RRj0Fs4
2CvyigLYuaz4mRXnllnA4DpbEn2mp5N5S0qHL3bC1ENRsOkcgm7Iho9xBhh7LVOW
/N/0cX5MO2R+AmoDTxQhVN5Xs93Zj6Xgn7rV3qn37D0G5qDGvoHuvz3P4foIolqW
1uicLZ47SA1Eqry/NkWsCKuMuR9IL7XGy8V9fmJ/mGyl/zBcni3VGkaVBEexEfoi
qKAe5HOaJNhGzFlZmV4MPxABAom+p6zJ7BtO1wXR6gUwfFMsCVqMrcWJqqYAxa/C
mpvoOur8UvgF3LyvXGmXQrmfdevF3psEhHFkh3ZupNND2SIBtY6bZuakke3gutr1
T7YQ8EG/S1VLHhp/TiYYHj/FiKhYKrvfIARBmJ5bYJ/mxrDmwZ2hYw8Q+TM92yjZ
f3h3xf+kxDQ5x/zLxK1eiyPxvflxT+CJAV2WBoQkefLDW8t5LR0HxCE52qfXFW5C
DKV2e3Wvwuit1eIJQs3EwqI9qYtMFhHJZlZ17EuQOBK0CjXDDYchOvZjZkB+UlK0
oDSdvVH4Ox/F999Ib+FoHysQUAIloLq8oYffNkHU2Ch1XzLIAIlfArFANR+wW20c
RB/O2j6PjrFLx3KhBkqdEBuZ2PckC1HnALcpiepDdEoxabRIW843ermXvK4d1JWJ
rmeawtyBKjhOc3wiQuHsVnI6UCrEWCHksC3nMT6jWjTp7+QxF9fP1uj5R6VbNZsE
VqQEtfPi7gTdHrdcDAMJuASBdE2qmHeF8jH6iKOXDp6TTKg/9TUX2u/KCPO5mWJS
IdlMG0cw9mIs7bz6z80AzeWI1zXqLWMryVT6Z+d9i9fmpDsEANCDgsG11iL531RU
aaglSQ6Q8H/9f1X2eHb7q1sj1couufDYBEwSBOB5YCdK/VUK1PXiYJBIE/voIx+B
aYJk8b8Yju/EjebY0JMjn1T4M7Mgf2BIHBXM6CNVRBToJPBpAcqiqzoJR1H6o1te
V6DKtKOGQmbzAtijo5vuRbu5hTxwYoALHEozOC/vucendm3i4GBXi8h5w+SpHFN5
qthSu1xPpOtbgsNdFdLbKsT5W5EHKB5zJ/GdWfO5I7ebZ61kDbZd7XJXkE3AUT2u
mOP5yKYxUofRyW863DBYTFDNG3awbsyVjn7lbKOVrzlUwHvNt0mPfJPkewmo5DpA
5gAXkfRqknNeJBO9IOWmcPdNjAj3P6LD1OR+bx8icLujUVD8ibwvPXYzRox9L5U6
ypQCCAyKBEqyVfD5TMRm+/Spx9tqShpll870mj73LQQYE7YSeothlPXd6Qomcf19
7dUtAtUbn/q/NbNQq6vOW3SumuM1We6X9FLua3EzNkxz8JZPRUbuvc1hj/HsSEBt
m4MoKj97H6Hx8pFVhz0CeqFllxGcsI1e4ySsZiVCRsDdenDBu7TQBS3T0DkS3l0W
wZ3U60eDVsiKnTOPNTnwVGDjFngOU8/IRu3VcpEmtiXxDbgOadt5birWdI2sEkPN
tbIR/dW+Vbi7sg7nMUWgqpYNUf2BeZqj4mkVjGu2GxvQUYlR5Db0IASxpdKyAC86
P66WYJZsOS7Qpt+go59hYy4OW633Ax2ARHJjkinuxCgIYMy5fszOEP6Ev9aa+c6j
stWnHTUIvEsfHsWZ27lt2S04SeIumMMNCFmnLcUzmPnOZ884xWuRa+iAzCbg7FgY
7WwGT16j5G3eHd23uda3QKAwCd/s3HfCrXdOIns3txRCRo2Ff1hYxkh3tRiwrjcG
bcGCiOUSMqoBHoTLkRaDa0S4L0KxJTsTdVlw7A+76oltBL+kRefR5SHYSiaULq3J
ou+N2Xe2QSMPbKePdd7erwPrGykFA9P+q4JMdEjvcBDgtBM0saYRgCitsstSbSuU
U6yeVvwd3k6S73eGyPH98O4VcF8NduNBPIhHDaGwKr1487F/crsmiaM133En/2md
mmKVHIGPHTmA1GOcQM3i/aLeW5GmnovmGL787WSaacW+1XLa0Eqn1+awlTJjsVPl
OrFvHdjmQVIiKdWfbQmkQtjXPZXLvKt8gVaIh14Uz6iLoAiO0Umpd06yBvfi1R0O
+dDb4QqHzTmBHlBL6VwwUBfo1WBbzRMXws4+nSrG13MTDO9fVWilS4imAMpJQ2dT
Dx2IBqXokcxCFw4EpBnXGi76myfzbKvov5nAw6HsSwUiOqv6dPpK03cE857ltmG5
H8Ckgr+A1bGkSTAIiNRwfGttYjcVJEzLSEJ0Ou//q+Oe7wwMeYkkFS8DXmZl1xab
Y8LK9SYM9fXXX8fv1ApLAmx7eqg6Z7jwEvCKKElAxcOI62rhVb9o9kuhIaIGgvPf
wabReaQvnoC6dESza8bbJtas0NoD9lH04TBQw/iPS8Pgk23CldmD9qqL3OWQOPmg
2NAd0m1yLWwH6ORRrNZaqA8n4IedMPwz2V57UxQv82u6dyvRytKkTuDYzXsybFe1
ZEsJbkhEvhJgTUNjKY4dKFrXftzGCaXBMrn2+T61j+teccy0m3WqQpe8L7MlUkQV
30vmF6S9UOm+EZ4BkUPQSLR+vio1PHbV0MnHrRrwnFlinMiXFSTAV+4fNJ1zNyBt
+pxa63YrUfTnEv7rpztAQ4HNHYUALfcOV6CW4IweeHYNdMZXDtTAdQZhKa2PTTfx
cMQXUcCoRTokMwnyI3qYh4M7Z32IILpvUTYuonWovyMmgSN5gVRYsF8cSyelxSKv
6v9rinHLsua7tThJehB4PNLbhiQxh/1JGYgOrCXGGLgeqgU6y/8LTaJ34UKzmHv6
DO0+UKgDHn699SGKzue6VvDTZG0gp9E9nlxZZfMWLGdDvS8SEqhlHLAARqt1g4ne
o098hNig0JmCYwtSwYg6Yuq+hu/oyf1YIQcwIw0+UchmgpPZ9M0EdR+1ahzclBfv
31uS/G5spUzS6tUoIqPJAliiG/eC4hLmOHLLWABpT97jsu/3s9eT1IAtQrxMWcUC
PvBS1v+dJkCPY7CqiPOAXsWuGXHznTRlJNBNOJH0uFRgO0EqgBnSVsOrArfvn2MY
usTMsvUbFZA6dLgUPfM/3KFRM247kvRlWtp3kmYcw6HPsSOSym9wI12ZsTdKHoWu
76DbxlIUIFjamHHedRQVzRFmjpjaaQJz64bsrGIAmqU9T4mv8nF1WwiQaS5cOa0h
PJPAosP4IJ5IJxh8xCeL307v8e4v78ETQqpx1bU5MRLPvah3CR3Huqt8xlQLzhPU
p9Afl8q7W3TiRjX7ePLz9ySSELXhXlvnjtPPn5XbsLYanurpB0vS4DaObWz2hkUH
4ij7soNEGDsZxIdHnQwl49g3NJ/FBJq01nD6cV6OdpK0E1JcnzqS4gab8Z+EHX7P
RCDCY07vZ+Xwjn18HXrzBw0yI8PFM2MzuxBQUO35v4iOuyfxxBVqnc8oHoACd1uu
EbXC2GpWhec4Ucs+kyX/Ysw0RsxPXXiwQIpTGjGvkRFHGvxSkb6h5gH3F3LZT3Sz
9ZShzb1+RZhQytwRomhLRgQULIQIxAy0L8EncgGR2mnRAylJmVGHIkj6050Cwprb
rWFCjUolsQ0VhVJyA0GVTeZK7hn+K33N0M8PzugfJpz1hwXGWppv5J2lU4jfAojk
KfQPSjHPmZNZemfE1aAXrmAUqrAtsyG3gHUJSrn2g7cJFzd9oCR/t3uBxmyvszZ6
LuM8rBmQMe9qvfFSs6/95nQXaj6tZCmzQCrUMdh/JPMxeoQ5x55l1qV1foiITLT+
9i0HncFS5NQMILm4Ye6u6+s3r5GysT+Dnw1NkmyfQUY+Kzm140ENoRNLLH87KCoO
5+DDG9ImUqRK8i2lqDcoPn9wc2UUiqNFk7K2fnroa88BfkLQ6wrsCNRRfVJO16G5
Bm8EXeLFCkb5P2m9ASJS4lodgsbUYsz/v1NiigTLoZaRehJD0/GWHyLWt9bfhhiS
nX/UBm7PCev7ycnzkF3Hdy1PUXsx16KB2jwCtV6dbldrMG7ltJw9/PGEXf9r8cAH
VWsPF+57OrSk3vsPJR6TccR2uTvLTO5usdVFH8Rjok3WGmM7ViA0P2CwXSBb7eoC
eTV3mrffLvA5lmCcTzU37p6VBDcdPxiLAUcdA5e7fU1r7EMlLSiax2jrJAwPysdh
CWQbLHYYuLRJ4yR89NrVBb2Z2BaD9UWGYh1GbvyMpgquPxUJXMPVkDbTB2Uzo11K
2OB/ECuPAhBJNJFgC4yTSEfiDPqNNKxyrLM54NHXVLmZO/a1pqqSTsuT8VCTBNNV
/4egj/SMgYGKj3q6UEYrqdX0Ky6yvk+y64GRD4fe5hNEHV1cZeLLx+2nRTBqxq5V
FcS193qrCnWukLXZJYSpc28ggYtwbwpp7cfsPM4lluRjDuavUruGh1tkoQt9T0Pz
SLANzGvekIwIrMuP4eHVm1GY7DkKiTCrEt9H+rsZ8cf9xJLgZYKG3Inbj5R/rFAi
HL8YjQyLXy6qvTQazrlPqSobuv5jb0VVQkyEDBAmRZZyJr5jwVpZJoIL69qDBDue
KO78SBge+wHKxZGYxGF6oBJw0YN/rrh3IKgjul+30yk/JLzzxCg1TDpNbb2P9DZm
1La4OmeoqJPKrrY0lrccQFR1sNikE+NisDOFv3JVP6t4he70em9n4FXhcje8KewA
P+6rLmpw92DLP+FuQ0Bd6Wq1MhX/TI6RtLavCsiKYgJw1LwtOvfYf/8cJ49cNK2W
HJpZCYKVNgvW8dT6zzckttA7pypb0SvnlgHZte2+U8mNLaAYKkk50geOFKottOhL
IysNH2iKeeF5JvQA9miclFPTjRc7ZdNyCKckGMqt9ZUc8ndN3f2epW4FgvlxyiUC
QtcD0QbNu+bZvsLeUpYSvCJ1RWAq/W+VkiCyZTyqCbnRkbbsPrwk9Rh8oUpmhZZj
Is7XEeU6Gar0T8c6pahj1MWL3fI4X7m08O3JOfcQDbPOIzrLjaSThyUOHFygF4lq
QpWQO9xuy/QNXce2rEPHu7yo7V4zvh3+M0Pl+9dr+Con8RLmnftgrPX1gzAryGST
jJoCSfrxn/Gi8rv3GCdXTiJ8QN5rQaMjRtJEa7jWeLLyrvzkyyh9BppV2/RX9mhz
MFj8djhOJJxJICLupTKP/C/liqLGP1MltGBn37IvXKLzBimg85uDCI1nf8cLPEQK
0a2df9OVsNqLfUJnFevHXl79L2tVlVEyVBanoUzWNjGoVgjyyp0K6Heub/3Odw+m
UF27IjjxRnX8kOG9bBqWtq58ERX1SD0NY9FMWHWP3+UU1Yus0C97QjRI0m28Hu3k
HKJwK5FNtyjXtwr8TTKJn5lRMS9SZih4NpIJ9kR7bNuJ7RMxbZr7ES/N44/HHOJU
QpFZHhZUrbqHBWEIDca6cb32uxVWrpHEt6jIaT2LgVTFnll9Vp8EXeSh7sbBzRxi
sw1DG1gt6sY8Y6f2LaqS90q8fFecVZ7x36lef1+n9fZKJuhwmqnHMGTVg0N/UHpU
azlbtIIqnJUaOSZvycE2+0aQbJ9umZe1upipyisIIfHer0BxcUagosfShV/2r/qE
tQ23CnlxiarnOnnOWETC7/AJFnjAjtpqkw6NTJSNUeOt/tPx7c2iA5QE/oQJ5hoB
4BhmopfD3eUudJql8dIWqh+dblMSfqTyaemd9UCb+FdP+UXlipGzcsq7kZG8qG97
njYM90us+jCyPUdCeaYhUYyNxyAWwOUl42SS5+WINOUq7Ic+Tv5fmIfymrbAsDE+
U2xZnNYMe1MZYoHej4bgUN9jTdm4ViZDfLMgHlsAna+Se2PVEL/XYVfP6yGH3sFQ
e5zrKyQeCWg/9kUjRzFGrp/8Ca8zPaLVwjq8ncQp2g8p3yRW3SzTRWCgmCqNz7HJ
FZxX8XV1y766zLkbznfYO3UMS+OvQOf5TSUTlHpCbBnlPYrnCvUY/alHmWt4E06R
AnIwvvDufbffamabzfZ9hf4sdA409eVa7UmnkCjDxDEYiTcnrGHkqOfOHlEWiwBh
Si+/acbLk5vdWIdcA6zX9oshEHHjYo5UlMrVcGsXDsvf/hsjDBVL1gvBRkCNTLx0
n6nVVvPrYDoZ/R6gO4cLGs0Cdz15jGzmTsP+Nn417/A4NBjXAKi3OLm5fPQxPFuO
OdwvoO6lcua3e3DMRIsT2J/2c4KKZ1nPKcwY5XHfBlkikgNGChE6U0QOF8LkJjHh
AUfX1J56GaofuMOgHGamDSPRvQ0tOYL/CBvoyB2cPFVImLH7fQFOXsn3mHxekCRp
GnJpj6DdISQSIGs5N6/q+nhCXzVwQ2tqV6vJddpr0u2pw9AhAUYIUGOWhoKBfYNy
BbJ4BTXMe7kTbH03aisINdvqPMwTrA5CZd0V9h8UXNDURgv72ID6DYjhWyKu1YxH
U4XVlm5uKwV9JWxbVN3Wf7fSjGPjSdc9t5sIJl34oLmWBLec66Zzc0+vdnlOhSuf
2oq8QdJFVJTd2I0ZkM/8PZ4aAB73L7nZjx5o12KnBbsa29h9Igtr1dUVcck+y6Mr
fgTsRHIJcaEN9jSOI4yksoQAlvdwiT0eD97J+MzgtPnKUr4dZwa+M9HKiCkWoyba
laKbMbU+id9GScPov71jg2CWBIk6xNyxvb5EzuhVxrGu0UYZgcAwuKqwZi5broK/
w/AIkv7LnrJnuOgCbp6Cm5fYmnxuHwRHwFNdikniHtf4HEpQKYvCyAFkbGijS5QV
P0+gIEYaPB5FUCe4mAticaab8Cv+qNT5aT5/YUdwS1jBqLyRYR48NqFNA4ccXHPS
iPYlPVsDlZ4K9roXukSyXTud+WQweEpYa7MR13uOnm6Op9fsu4DIcTNtUdv78ihq
tzQimAJbFI+hqR87N+k4r+LIuq/G8QuwFyVl9G0qKH1SwZMGaK8pNMlY6/mBnJbi
gAmqu17f7hri+gIzJPyJd/0BPKrh/OWLBHbJoRCIQ/Cu/sy/W3KkYjNDqw5WwjNy
qGRtaIY2u/CTSWnIc+1PF2WC4KXmo9oz/CLr/65EIs+j2IDLJchxN7JnRkaOjz0W
CoyG74gUHNPfsiVamjt5wUih9cuxdlr+ci0GcEPXIR10Fb91Fna0uMOFjvFhxp1g
T6JRRjieKUYucbSy6KazyJSGfZnzDtitJ5KYIf9EvDrfeCygwSccNLuu9UMw0n5i
QYvC2DGSqLqlLo7htzA0BI5vABmWZilK45JdAPoq0eJkSF12o7vmHLf6/MSyS7hR
hJev9CXb39+J6PW9+f3ZpHtB9jSmNygynDiWOlOPqa2t2kiaMPSegTj7dxGwPjB3
JekMwinZf4e/HBUFw+2D082pfdhKn7Zvr24XbJRxA78EDUsbNWiY1px5Ji8HWyke
dA7rvAb3UFleFaSdI9YKwABkara00KQYYQoA3tuNwuT2rqCEWxhmc8vdqPRgX8CB
so3Y0XsaWaWB0H349jjTJhjF7mJgaOWLlhV/dcsuo5zl7LS8BQujh2z4TF3yrtgV
vCt6FQNWP66M8N9h5mOIF2O36R78gZGA8Y4XZaG6qcAJ1GkyeFwwqYU+qriEe+D3
iXzZez35/K89a67vRRBSijDes+kjPhulUzgSCCBpN6Nhc/izgpp59wXWAoQ9/UlZ
agTzURZD/8i6/xUyV0L0rdunLH5DVkRJcCVY2kRHNQ9vCb5l6DFmYn7ETxHzFbUq
5iI4EKJ1hYO59zvA2bXwmh80F9d/bmk2qejXayNYMiV+vAsjzbDc4YekirFTM55n
lUrRfYAF5Vx5kYchzEjgVnQPQtljV7S5Y4AvhB7vihepEhCh3onDgzwLP77O6swQ
KO7wbAiLWK3YhMnzHF93SNXbi1k7yx3Frlu5c1+M9dhAvxAH917Y2djMP1s5R0Ny
k0z+AP24p4IrTu6jl7LiwCsMa5sMm5TYPiABSAdFE4awbAaRmSSFiJr+qyWct4KV
EXlRD9lgZzTL5EbXs/0ZrFwCW+MVM+o5g1RhJuBFTgKi+cmyBLKAxUZSZ+IQMmD1
0QNGc9Uivc6+KvuJH59r33RK2nI2qC4o1erOz4vS5REz5r+yJ8s9/P0ehA9aRmwL
Excyn2v0JJD9qDT8SIWW6nl7cP66+tqX5IXXlnsbTfiPmXVCK6VcMfhUVKvZD8ZA
ykN5qmiL/LmqL8HgLDcqLs6y1VNqT4eMo2YJlE/f7dzAVWVsp4x7zOVe1L2y0oBh
hfPzOLQWNYrIMJHMcLhGPaEJooMATmpsLgdEPexlKqQOZNGsFDOURKcG2qHGus9j
tu3UMFUijUVKLMyXz6W/DKg4ZrC6VH4KOiRwQItxR1brPkzGKKh5iGZnJASFICsq
2aGxeq9XVsWtEPlI/xwUfZ++tyPDUW7QYabpQSqNRUcGLo3pL41X9x1SxuKRFpe8
2BxE4EwoH8yj5LqN44RuQQTFO/poDKLSj0YMyyP6+H97i8PWPfxzw8FC15ZgEVw2
GhsjaMH5Bx7L8BiUC6xIQydwfGhbD7Pou1nkxWwr5fl47EfL87aMsYdsciuWBfHE
Xr0QqurjN4HQi6l6LSoOPTM0JvHH4nirru5oWIZAo0RKOdEjdo1WfjGTXCzkN/DM
j6qcYaH5Cf99xQn03tmYRmDxzbTm5H6tgYJyCY7Tacj+6Fw9MXPW7rZK9LJ+e/eE
zawKGrJKRx226cy8ye+1sNThHLHXjIKm721KyRNH4xovvIwGG5aWBc0heQ291+q/
sc3lwY9SBxYw6vkYtwi8lm41WCayrUORgHDjF5ZV2lZT0lfig71F10FnZ6CnutEs
2eWfy8PnmWUphS1IBk7nZoEWoJqODBYyD9fvlQAoeItIeQ+mCn7GFJw02BK+5N2u
zNf9CEtnUgD1GUTf+IGJHjWd0HLSo9EwiB7IFg/cG27Rke6qC6COGWztVeqMIP4m
3uvt1uZpXOLrTK3HDNVfp+iEoliIl20iq/kLQXZ39oYHY01klWKe7Jzqx0QGGEcV
/Fr9DIGz4lP1w9Tvi5QIdPNR51ajlrjge/8ZfD8rlbWdpMW0AzdcdsCM8x1dwHTR
65PstE0DGuspbBZK4ll32Sh6yVVFE13vE+GU3uULg6e8CLv6yYY+wSf/l+kSKZgF
+8mQ4scX4s0a9KtTouWreJme5XPFxWbM6NRQRSKzBj3ZizqHg+MkuzOxVY+VbDiY
eBUawtw2h8UZc0iglcIVqY01f+pQbp2kilaFGxEu4dpwv1PLPEJMML8klP5v0Spd
HpygOyLybDEbzAR8/v8GF9pBf/EeVtGLT9SjjMM3cIxvnoCF0n9BVB0ZkqOl5/tq
FtGGP2LTZ88f4MRO/t6g54jjNrtMf3Ju4rQkdplQDXZyIlaGpDT47UBEF84ED0EO
PlHcFBaWA+d64sgvzrmDZe1yLmUpWrU5drqpIoRm52gUgbX2oJCX7QnKSNJCuLk1
3SlUsB7g2386k9CSBRFur0bSR1mHQ8k/e67CYXXPA3zhvmI7YBJogEEqqLdTcWca
2+Hpvzln6ts9SHPw27pezcoF6PSkdoMnKmCrJkGmdwLE+dgPURhF+N3Y0PL2p4z7
rG9v5y1BRCpEIZIX3e3N/GuYzFJezOt23508UeBvyy+ZT++fnnc1LKdn48oZ05on
YZUO2xjhddxIwstqR4RdJ9khCWhNEMr+h2HP45zXLeovz78Kwf93YgmYah/XDc2u
tz9OCCDOfd3z5x0wy4S+LLcPU3HLKexlHAyJcMr6oPfh0IWBN9D5HK5ieysNvdPr
JZoDgwRpZx4aPLvChJAeB9GRoZ+hBx3nIFU4DaA9NZrJ3T59XEAWydoCZMAvvx+F
hmv0pVzodE3GyuQj4NE9RHBw0lM2obqRhD4WxHnPii22hxQ24X47OtWy+asLMjte
6apRrSqKkpg2nnPi6ZrNlu44N2XyVE7PEaC+qVYJTdRoDJUtI1PaOMYiOdG2RL/+
rYYQBMwvDS1TehECjL79mK1cRrl/pNYFfUp6aKGKK3Xu5ankOyno2yh3HX+bhB9/
WOlrEHZfQloiZs9CZdISk4AVpQzb7wfQzTd/5WiUeDeojxZDlHYITTQJTouObHdE
TIWbf9D8xs7m04wlrZY5HX3Gd5OpxDgO3XYX0Vy/kxc=
`protect END_PROTECTED
